package enc_8b10b_pkg;

  // MSB -> LSB
  // typedef struct packed {
  //   logic ctrl_symb;
  //   logic disp_front;
  //   logic code_err;
  //   logic disp_end;
  //   logic [9:0] symb;
  // } enc_symb_t;























































































  logic [13:0] enc_symb [0:1023] = '{
    // ctrl_symb  disp_front  code_err  disp_end  symb
      {1'b0,      1'b0,       1'b0,     1'b0,     10'b0010_111001}, // D.00.0, disp_front = 0, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b0,     10'b0010_101110}, // D.01.0, disp_front = 0, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b0,     10'b0010_101101}, // D.02.0, disp_front = 0, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b1,     10'b1101_100011}, // D.03.0, disp_front = 0, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b0,     10'b0010_101011}, // D.04.0, disp_front = 0, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b1,     10'b1101_100101}, // D.05.0, disp_front = 0, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b1,     10'b1101_100110}, // D.06.0, disp_front = 0, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b1,     10'b1101_000111}, // D.07.0, disp_front = 0, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b0,     10'b0010_100111}, // D.08.0, disp_front = 0, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b1,     10'b1101_101001}, // D.09.0, disp_front = 0, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b1,     10'b1101_101010}, // D.10.0, disp_front = 0, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b1,     10'b1101_001011}, // D.11.0, disp_front = 0, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b1,     10'b1101_101100}, // D.12.0, disp_front = 0, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b1,     10'b1101_001101}, // D.13.0, disp_front = 0, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b1,     10'b1101_001110}, // D.14.0, disp_front = 0, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b0,     10'b0010_111010}, // D.15.0, disp_front = 0, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b0,     10'b0010_110110}, // D.16.0, disp_front = 0, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b1,     10'b1101_110001}, // D.17.0, disp_front = 0, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b1,     10'b1101_110010}, // D.18.0, disp_front = 0, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b1,     10'b1101_010011}, // D.19.0, disp_front = 0, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b1,     10'b1101_110100}, // D.20.0, disp_front = 0, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b1,     10'b1101_010101}, // D.21.0, disp_front = 0, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b1,     10'b1101_010110}, // D.22.0, disp_front = 0, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b0,     10'b0010_010111}, // D.23.0, disp_front = 0, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b0,     10'b0010_110011}, // D.24.0, disp_front = 0, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b1,     10'b1101_011001}, // D.25.0, disp_front = 0, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b1,     10'b1101_011010}, // D.26.0, disp_front = 0, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b0,     10'b0010_011011}, // D.27.0, disp_front = 0, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b1,     10'b1101_011100}, // D.28.0, disp_front = 0, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b0,     10'b0010_011101}, // D.29.0, disp_front = 0, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b0,     10'b0010_011110}, // D.30.0, disp_front = 0, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b0,     10'b0010_110101}, // D.31.0, disp_front = 0, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b1,     10'b1001_111001}, // D.00.1, disp_front = 0, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b1,     10'b1001_101110}, // D.01.1, disp_front = 0, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b1,     10'b1001_101101}, // D.02.1, disp_front = 0, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b0,     10'b1001_100011}, // D.03.1, disp_front = 0, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b1,     10'b1001_101011}, // D.04.1, disp_front = 0, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b0,     10'b1001_100101}, // D.05.1, disp_front = 0, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b0,     10'b1001_100110}, // D.06.1, disp_front = 0, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b0,     10'b1001_000111}, // D.07.1, disp_front = 0, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b1,     10'b1001_100111}, // D.08.1, disp_front = 0, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b0,     10'b1001_101001}, // D.09.1, disp_front = 0, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b0,     10'b1001_101010}, // D.10.1, disp_front = 0, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b0,     10'b1001_001011}, // D.11.1, disp_front = 0, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b0,     10'b1001_101100}, // D.12.1, disp_front = 0, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b0,     10'b1001_001101}, // D.13.1, disp_front = 0, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b0,     10'b1001_001110}, // D.14.1, disp_front = 0, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b1,     10'b1001_111010}, // D.15.1, disp_front = 0, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b1,     10'b1001_110110}, // D.16.1, disp_front = 0, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b0,     10'b1001_110001}, // D.17.1, disp_front = 0, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b0,     10'b1001_110010}, // D.18.1, disp_front = 0, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b0,     10'b1001_010011}, // D.19.1, disp_front = 0, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b0,     10'b1001_110100}, // D.20.1, disp_front = 0, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b0,     10'b1001_010101}, // D.21.1, disp_front = 0, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b0,     10'b1001_010110}, // D.22.1, disp_front = 0, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b1,     10'b1001_010111}, // D.23.1, disp_front = 0, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b1,     10'b1001_110011}, // D.24.1, disp_front = 0, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b0,     10'b1001_011001}, // D.25.1, disp_front = 0, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b0,     10'b1001_011010}, // D.26.1, disp_front = 0, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b1,     10'b1001_011011}, // D.27.1, disp_front = 0, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b0,     10'b1001_011100}, // D.28.1, disp_front = 0, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b1,     10'b1001_011101}, // D.29.1, disp_front = 0, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b1,     10'b1001_011110}, // D.30.1, disp_front = 0, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b1,     10'b1001_110101}, // D.31.1, disp_front = 0, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b1,     10'b1010_111001}, // D.00.2, disp_front = 0, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b1,     10'b1010_101110}, // D.01.2, disp_front = 0, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b1,     10'b1010_101101}, // D.02.2, disp_front = 0, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b0,     10'b1010_100011}, // D.03.2, disp_front = 0, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b1,     10'b1010_101011}, // D.04.2, disp_front = 0, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b0,     10'b1010_100101}, // D.05.2, disp_front = 0, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b0,     10'b1010_100110}, // D.06.2, disp_front = 0, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b0,     10'b1010_000111}, // D.07.2, disp_front = 0, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b1,     10'b1010_100111}, // D.08.2, disp_front = 0, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b0,     10'b1010_101001}, // D.09.2, disp_front = 0, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b0,     10'b1010_101010}, // D.10.2, disp_front = 0, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b0,     10'b1010_001011}, // D.11.2, disp_front = 0, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b0,     10'b1010_101100}, // D.12.2, disp_front = 0, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b0,     10'b1010_001101}, // D.13.2, disp_front = 0, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b0,     10'b1010_001110}, // D.14.2, disp_front = 0, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b1,     10'b1010_111010}, // D.15.2, disp_front = 0, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b1,     10'b1010_110110}, // D.16.2, disp_front = 0, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b0,     10'b1010_110001}, // D.17.2, disp_front = 0, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b0,     10'b1010_110010}, // D.18.2, disp_front = 0, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b0,     10'b1010_010011}, // D.19.2, disp_front = 0, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b0,     10'b1010_110100}, // D.20.2, disp_front = 0, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b0,     10'b1010_010101}, // D.21.2, disp_front = 0, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b0,     10'b1010_010110}, // D.22.2, disp_front = 0, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b1,     10'b1010_010111}, // D.23.2, disp_front = 0, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b1,     10'b1010_110011}, // D.24.2, disp_front = 0, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b0,     10'b1010_011001}, // D.25.2, disp_front = 0, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b0,     10'b1010_011010}, // D.26.2, disp_front = 0, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b1,     10'b1010_011011}, // D.27.2, disp_front = 0, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b0,     10'b1010_011100}, // D.28.2, disp_front = 0, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b1,     10'b1010_011101}, // D.29.2, disp_front = 0, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b1,     10'b1010_011110}, // D.30.2, disp_front = 0, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b1,     10'b1010_110101}, // D.31.2, disp_front = 0, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b1,     10'b1100_111001}, // D.00.3, disp_front = 0, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b1,     10'b1100_101110}, // D.01.3, disp_front = 0, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b1,     10'b1100_101101}, // D.02.3, disp_front = 0, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b0,     10'b0011_100011}, // D.03.3, disp_front = 0, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b1,     10'b1100_101011}, // D.04.3, disp_front = 0, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b0,     10'b0011_100101}, // D.05.3, disp_front = 0, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b0,     10'b0011_100110}, // D.06.3, disp_front = 0, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b0,     10'b0011_000111}, // D.07.3, disp_front = 0, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b1,     10'b1100_100111}, // D.08.3, disp_front = 0, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b0,     10'b0011_101001}, // D.09.3, disp_front = 0, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b0,     10'b0011_101010}, // D.10.3, disp_front = 0, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b0,     10'b0011_001011}, // D.11.3, disp_front = 0, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b0,     10'b0011_101100}, // D.12.3, disp_front = 0, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b0,     10'b0011_001101}, // D.13.3, disp_front = 0, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b0,     10'b0011_001110}, // D.14.3, disp_front = 0, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b1,     10'b1100_111010}, // D.15.3, disp_front = 0, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b1,     10'b1100_110110}, // D.16.3, disp_front = 0, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b0,     10'b0011_110001}, // D.17.3, disp_front = 0, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b0,     10'b0011_110010}, // D.18.3, disp_front = 0, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b0,     10'b0011_010011}, // D.19.3, disp_front = 0, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b0,     10'b0011_110100}, // D.20.3, disp_front = 0, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b0,     10'b0011_010101}, // D.21.3, disp_front = 0, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b0,     10'b0011_010110}, // D.22.3, disp_front = 0, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b1,     10'b1100_010111}, // D.23.3, disp_front = 0, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b1,     10'b1100_110011}, // D.24.3, disp_front = 0, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b0,     10'b0011_011001}, // D.25.3, disp_front = 0, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b0,     10'b0011_011010}, // D.26.3, disp_front = 0, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b1,     10'b1100_011011}, // D.27.3, disp_front = 0, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b0,     10'b0011_011100}, // D.28.3, disp_front = 0, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b1,     10'b1100_011101}, // D.29.3, disp_front = 0, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b1,     10'b1100_011110}, // D.30.3, disp_front = 0, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b1,     10'b1100_110101}, // D.31.3, disp_front = 0, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b0,     10'b0100_111001}, // D.00.4, disp_front = 0, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b0,     10'b0100_101110}, // D.01.4, disp_front = 0, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b0,     10'b0100_101101}, // D.02.4, disp_front = 0, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b1,     10'b1011_100011}, // D.03.4, disp_front = 0, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b0,     10'b0100_101011}, // D.04.4, disp_front = 0, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b1,     10'b1011_100101}, // D.05.4, disp_front = 0, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b1,     10'b1011_100110}, // D.06.4, disp_front = 0, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b1,     10'b1011_000111}, // D.07.4, disp_front = 0, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b0,     10'b0100_100111}, // D.08.4, disp_front = 0, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b1,     10'b1011_101001}, // D.09.4, disp_front = 0, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b1,     10'b1011_101010}, // D.10.4, disp_front = 0, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b1,     10'b1011_001011}, // D.11.4, disp_front = 0, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b1,     10'b1011_101100}, // D.12.4, disp_front = 0, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b1,     10'b1011_001101}, // D.13.4, disp_front = 0, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b1,     10'b1011_001110}, // D.14.4, disp_front = 0, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b0,     10'b0100_111010}, // D.15.4, disp_front = 0, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b0,     10'b0100_110110}, // D.16.4, disp_front = 0, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b1,     10'b1011_110001}, // D.17.4, disp_front = 0, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b1,     10'b1011_110010}, // D.18.4, disp_front = 0, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b1,     10'b1011_010011}, // D.19.4, disp_front = 0, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b1,     10'b1011_110100}, // D.20.4, disp_front = 0, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b1,     10'b1011_010101}, // D.21.4, disp_front = 0, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b1,     10'b1011_010110}, // D.22.4, disp_front = 0, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b0,     10'b0100_010111}, // D.23.4, disp_front = 0, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b0,     10'b0100_110011}, // D.24.4, disp_front = 0, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b1,     10'b1011_011001}, // D.25.4, disp_front = 0, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b1,     10'b1011_011010}, // D.26.4, disp_front = 0, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b0,     10'b0100_011011}, // D.27.4, disp_front = 0, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b1,     10'b1011_011100}, // D.28.4, disp_front = 0, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b0,     10'b0100_011101}, // D.29.4, disp_front = 0, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b0,     10'b0100_011110}, // D.30.4, disp_front = 0, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b0,     10'b0100_110101}, // D.31.4, disp_front = 0, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b1,     10'b0101_111001}, // D.00.5, disp_front = 0, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b1,     10'b0101_101110}, // D.01.5, disp_front = 0, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b1,     10'b0101_101101}, // D.02.5, disp_front = 0, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b0,     10'b0101_100011}, // D.03.5, disp_front = 0, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b1,     10'b0101_101011}, // D.04.5, disp_front = 0, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b0,     10'b0101_100101}, // D.05.5, disp_front = 0, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b0,     10'b0101_100110}, // D.06.5, disp_front = 0, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b0,     10'b0101_000111}, // D.07.5, disp_front = 0, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b1,     10'b0101_100111}, // D.08.5, disp_front = 0, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b0,     10'b0101_101001}, // D.09.5, disp_front = 0, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b0,     10'b0101_101010}, // D.10.5, disp_front = 0, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b0,     10'b0101_001011}, // D.11.5, disp_front = 0, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b0,     10'b0101_101100}, // D.12.5, disp_front = 0, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b0,     10'b0101_001101}, // D.13.5, disp_front = 0, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b0,     10'b0101_001110}, // D.14.5, disp_front = 0, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b1,     10'b0101_111010}, // D.15.5, disp_front = 0, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b1,     10'b0101_110110}, // D.16.5, disp_front = 0, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b0,     10'b0101_110001}, // D.17.5, disp_front = 0, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b0,     10'b0101_110010}, // D.18.5, disp_front = 0, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b0,     10'b0101_010011}, // D.19.5, disp_front = 0, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b0,     10'b0101_110100}, // D.20.5, disp_front = 0, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b0,     10'b0101_010101}, // D.21.5, disp_front = 0, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b0,     10'b0101_010110}, // D.22.5, disp_front = 0, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b1,     10'b0101_010111}, // D.23.5, disp_front = 0, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b1,     10'b0101_110011}, // D.24.5, disp_front = 0, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b0,     10'b0101_011001}, // D.25.5, disp_front = 0, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b0,     10'b0101_011010}, // D.26.5, disp_front = 0, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b1,     10'b0101_011011}, // D.27.5, disp_front = 0, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b0,     10'b0101_011100}, // D.28.5, disp_front = 0, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b1,     10'b0101_011101}, // D.29.5, disp_front = 0, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b1,     10'b0101_011110}, // D.30.5, disp_front = 0, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b1,     10'b0101_110101}, // D.31.5, disp_front = 0, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b1,     10'b0110_111001}, // D.00.6, disp_front = 0, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b1,     10'b0110_101110}, // D.01.6, disp_front = 0, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b1,     10'b0110_101101}, // D.02.6, disp_front = 0, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b0,     10'b0110_100011}, // D.03.6, disp_front = 0, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b1,     10'b0110_101011}, // D.04.6, disp_front = 0, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b0,     10'b0110_100101}, // D.05.6, disp_front = 0, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b0,     10'b0110_100110}, // D.06.6, disp_front = 0, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b0,     10'b0110_000111}, // D.07.6, disp_front = 0, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b1,     10'b0110_100111}, // D.08.6, disp_front = 0, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b0,     10'b0110_101001}, // D.09.6, disp_front = 0, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b0,     10'b0110_101010}, // D.10.6, disp_front = 0, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b0,     10'b0110_001011}, // D.11.6, disp_front = 0, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b0,     10'b0110_101100}, // D.12.6, disp_front = 0, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b0,     10'b0110_001101}, // D.13.6, disp_front = 0, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b0,     10'b0110_001110}, // D.14.6, disp_front = 0, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b1,     10'b0110_111010}, // D.15.6, disp_front = 0, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b1,     10'b0110_110110}, // D.16.6, disp_front = 0, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b0,     10'b0110_110001}, // D.17.6, disp_front = 0, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b0,     10'b0110_110010}, // D.18.6, disp_front = 0, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b0,     10'b0110_010011}, // D.19.6, disp_front = 0, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b0,     10'b0110_110100}, // D.20.6, disp_front = 0, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b0,     10'b0110_010101}, // D.21.6, disp_front = 0, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b0,     10'b0110_010110}, // D.22.6, disp_front = 0, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b1,     10'b0110_010111}, // D.23.6, disp_front = 0, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b1,     10'b0110_110011}, // D.24.6, disp_front = 0, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b0,     10'b0110_011001}, // D.25.6, disp_front = 0, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b0,     10'b0110_011010}, // D.26.6, disp_front = 0, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b1,     10'b0110_011011}, // D.27.6, disp_front = 0, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b0,     10'b0110_011100}, // D.28.6, disp_front = 0, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b1,     10'b0110_011101}, // D.29.6, disp_front = 0, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b1,     10'b0110_011110}, // D.30.6, disp_front = 0, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b1,     10'b0110_110101}, // D.31.6, disp_front = 0, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b0,     10'b1000_111001}, // D.00.7, disp_front = 0, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b0,     10'b1000_101110}, // D.01.7, disp_front = 0, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b0,     10'b1000_101101}, // D.02.7, disp_front = 0, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b1,     10'b0111_100011}, // D.03.7, disp_front = 0, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b0,     10'b1000_101011}, // D.04.7, disp_front = 0, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b1,     10'b0111_100101}, // D.05.7, disp_front = 0, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b1,     10'b0111_100110}, // D.06.7, disp_front = 0, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b1,     10'b0111_000111}, // D.07.7, disp_front = 0, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b0,     10'b1000_100111}, // D.08.7, disp_front = 0, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b1,     10'b0111_101001}, // D.09.7, disp_front = 0, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b1,     10'b0111_101010}, // D.10.7, disp_front = 0, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b1,     10'b0111_001011}, // D.11.7, disp_front = 0, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b1,     10'b0111_101100}, // D.12.7, disp_front = 0, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b1,     10'b0111_001101}, // D.13.7, disp_front = 0, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b1,     10'b0111_001110}, // D.14.7, disp_front = 0, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b0,     10'b1000_111010}, // D.15.7, disp_front = 0, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b0,     10'b1000_110110}, // D.16.7, disp_front = 0, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b1,     10'b1110_110001}, // D.17.7, disp_front = 0, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b1,     10'b1110_110010}, // D.18.7, disp_front = 0, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b1,     10'b0111_010011}, // D.19.7, disp_front = 0, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b1,     10'b1110_110100}, // D.20.7, disp_front = 0, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b1,     10'b0111_010101}, // D.21.7, disp_front = 0, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b1,     10'b0111_010110}, // D.22.7, disp_front = 0, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b0,     10'b1000_010111}, // D.23.7, disp_front = 0, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b0,     10'b1000_110011}, // D.24.7, disp_front = 0, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b1,     10'b0111_011001}, // D.25.7, disp_front = 0, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b1,     10'b0111_011010}, // D.26.7, disp_front = 0, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b0,     10'b1000_011011}, // D.27.7, disp_front = 0, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b1,     10'b0111_011100}, // D.28.7, disp_front = 0, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b0,     10'b1000_011101}, // D.29.7, disp_front = 0, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b0,     10'b1000_011110}, // D.30.7, disp_front = 0, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b0,       1'b0,     1'b0,     10'b1000_110101}, // D.31.7, disp_front = 0, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b1,     10'b1101_000110}, // D.00.0, disp_front = 1, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b1,     10'b1101_010001}, // D.01.0, disp_front = 1, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b1,     10'b1101_010010}, // D.02.0, disp_front = 1, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b0,     10'b0010_100011}, // D.03.0, disp_front = 1, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b1,     10'b1101_010100}, // D.04.0, disp_front = 1, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b0,     10'b0010_100101}, // D.05.0, disp_front = 1, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b0,     10'b0010_100110}, // D.06.0, disp_front = 1, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b0,     10'b0010_111000}, // D.07.0, disp_front = 1, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b1,     10'b1101_011000}, // D.08.0, disp_front = 1, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b0,     10'b0010_101001}, // D.09.0, disp_front = 1, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b0,     10'b0010_101010}, // D.10.0, disp_front = 1, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b0,     10'b0010_001011}, // D.11.0, disp_front = 1, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b0,     10'b0010_101100}, // D.12.0, disp_front = 1, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b0,     10'b0010_001101}, // D.13.0, disp_front = 1, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b0,     10'b0010_001110}, // D.14.0, disp_front = 1, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b1,     10'b1101_000101}, // D.15.0, disp_front = 1, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b1,     10'b1101_001001}, // D.16.0, disp_front = 1, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b0,     10'b0010_110001}, // D.17.0, disp_front = 1, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b0,     10'b0010_110010}, // D.18.0, disp_front = 1, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b0,     10'b0010_010011}, // D.19.0, disp_front = 1, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b0,     10'b0010_110100}, // D.20.0, disp_front = 1, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b0,     10'b0010_010101}, // D.21.0, disp_front = 1, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b0,     10'b0010_010110}, // D.22.0, disp_front = 1, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b1,     10'b1101_101000}, // D.23.0, disp_front = 1, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b1,     10'b1101_001100}, // D.24.0, disp_front = 1, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b0,     10'b0010_011001}, // D.25.0, disp_front = 1, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b0,     10'b0010_011010}, // D.26.0, disp_front = 1, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b1,     10'b1101_100100}, // D.27.0, disp_front = 1, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b0,     10'b0010_011100}, // D.28.0, disp_front = 1, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b1,     10'b1101_100010}, // D.29.0, disp_front = 1, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b1,     10'b1101_100001}, // D.30.0, disp_front = 1, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b1,     10'b1101_001010}, // D.31.0, disp_front = 1, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b0,     10'b1001_000110}, // D.00.1, disp_front = 1, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b0,     10'b1001_010001}, // D.01.1, disp_front = 1, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b0,     10'b1001_010010}, // D.02.1, disp_front = 1, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b1,     10'b1001_100011}, // D.03.1, disp_front = 1, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b0,     10'b1001_010100}, // D.04.1, disp_front = 1, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b1,     10'b1001_100101}, // D.05.1, disp_front = 1, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b1,     10'b1001_100110}, // D.06.1, disp_front = 1, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b1,     10'b1001_111000}, // D.07.1, disp_front = 1, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b0,     10'b1001_011000}, // D.08.1, disp_front = 1, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b1,     10'b1001_101001}, // D.09.1, disp_front = 1, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b1,     10'b1001_101010}, // D.10.1, disp_front = 1, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b1,     10'b1001_001011}, // D.11.1, disp_front = 1, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b1,     10'b1001_101100}, // D.12.1, disp_front = 1, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b1,     10'b1001_001101}, // D.13.1, disp_front = 1, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b1,     10'b1001_001110}, // D.14.1, disp_front = 1, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b0,     10'b1001_000101}, // D.15.1, disp_front = 1, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b0,     10'b1001_001001}, // D.16.1, disp_front = 1, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b1,     10'b1001_110001}, // D.17.1, disp_front = 1, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b1,     10'b1001_110010}, // D.18.1, disp_front = 1, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b1,     10'b1001_010011}, // D.19.1, disp_front = 1, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b1,     10'b1001_110100}, // D.20.1, disp_front = 1, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b1,     10'b1001_010101}, // D.21.1, disp_front = 1, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b1,     10'b1001_010110}, // D.22.1, disp_front = 1, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b0,     10'b1001_101000}, // D.23.1, disp_front = 1, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b0,     10'b1001_001100}, // D.24.1, disp_front = 1, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b1,     10'b1001_011001}, // D.25.1, disp_front = 1, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b1,     10'b1001_011010}, // D.26.1, disp_front = 1, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b0,     10'b1001_100100}, // D.27.1, disp_front = 1, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b1,     10'b1001_011100}, // D.28.1, disp_front = 1, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b0,     10'b1001_100010}, // D.29.1, disp_front = 1, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b0,     10'b1001_100001}, // D.30.1, disp_front = 1, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b0,     10'b1001_001010}, // D.31.1, disp_front = 1, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b0,     10'b1010_000110}, // D.00.2, disp_front = 1, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b0,     10'b1010_010001}, // D.01.2, disp_front = 1, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b0,     10'b1010_010010}, // D.02.2, disp_front = 1, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b1,     10'b1010_100011}, // D.03.2, disp_front = 1, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b0,     10'b1010_010100}, // D.04.2, disp_front = 1, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b1,     10'b1010_100101}, // D.05.2, disp_front = 1, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b1,     10'b1010_100110}, // D.06.2, disp_front = 1, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b1,     10'b1010_111000}, // D.07.2, disp_front = 1, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b0,     10'b1010_011000}, // D.08.2, disp_front = 1, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b1,     10'b1010_101001}, // D.09.2, disp_front = 1, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b1,     10'b1010_101010}, // D.10.2, disp_front = 1, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b1,     10'b1010_001011}, // D.11.2, disp_front = 1, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b1,     10'b1010_101100}, // D.12.2, disp_front = 1, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b1,     10'b1010_001101}, // D.13.2, disp_front = 1, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b1,     10'b1010_001110}, // D.14.2, disp_front = 1, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b0,     10'b1010_000101}, // D.15.2, disp_front = 1, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b0,     10'b1010_001001}, // D.16.2, disp_front = 1, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b1,     10'b1010_110001}, // D.17.2, disp_front = 1, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b1,     10'b1010_110010}, // D.18.2, disp_front = 1, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b1,     10'b1010_010011}, // D.19.2, disp_front = 1, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b1,     10'b1010_110100}, // D.20.2, disp_front = 1, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b1,     10'b1010_010101}, // D.21.2, disp_front = 1, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b1,     10'b1010_010110}, // D.22.2, disp_front = 1, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b0,     10'b1010_101000}, // D.23.2, disp_front = 1, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b0,     10'b1010_001100}, // D.24.2, disp_front = 1, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b1,     10'b1010_011001}, // D.25.2, disp_front = 1, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b1,     10'b1010_011010}, // D.26.2, disp_front = 1, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b0,     10'b1010_100100}, // D.27.2, disp_front = 1, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b1,     10'b1010_011100}, // D.28.2, disp_front = 1, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b0,     10'b1010_100010}, // D.29.2, disp_front = 1, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b0,     10'b1010_100001}, // D.30.2, disp_front = 1, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b0,     10'b1010_001010}, // D.31.2, disp_front = 1, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b0,     10'b0011_000110}, // D.00.3, disp_front = 1, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b0,     10'b0011_010001}, // D.01.3, disp_front = 1, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b0,     10'b0011_010010}, // D.02.3, disp_front = 1, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b1,     10'b1100_100011}, // D.03.3, disp_front = 1, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b0,     10'b0011_010100}, // D.04.3, disp_front = 1, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b1,     10'b1100_100101}, // D.05.3, disp_front = 1, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b1,     10'b1100_100110}, // D.06.3, disp_front = 1, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b1,     10'b1100_111000}, // D.07.3, disp_front = 1, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b0,     10'b0011_011000}, // D.08.3, disp_front = 1, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b1,     10'b1100_101001}, // D.09.3, disp_front = 1, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b1,     10'b1100_101010}, // D.10.3, disp_front = 1, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b1,     10'b1100_001011}, // D.11.3, disp_front = 1, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b1,     10'b1100_101100}, // D.12.3, disp_front = 1, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b1,     10'b1100_001101}, // D.13.3, disp_front = 1, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b1,     10'b1100_001110}, // D.14.3, disp_front = 1, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b0,     10'b0011_000101}, // D.15.3, disp_front = 1, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b0,     10'b0011_001001}, // D.16.3, disp_front = 1, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b1,     10'b1100_110001}, // D.17.3, disp_front = 1, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b1,     10'b1100_110010}, // D.18.3, disp_front = 1, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b1,     10'b1100_010011}, // D.19.3, disp_front = 1, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b1,     10'b1100_110100}, // D.20.3, disp_front = 1, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b1,     10'b1100_010101}, // D.21.3, disp_front = 1, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b1,     10'b1100_010110}, // D.22.3, disp_front = 1, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b0,     10'b0011_101000}, // D.23.3, disp_front = 1, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b0,     10'b0011_001100}, // D.24.3, disp_front = 1, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b1,     10'b1100_011001}, // D.25.3, disp_front = 1, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b1,     10'b1100_011010}, // D.26.3, disp_front = 1, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b0,     10'b0011_100100}, // D.27.3, disp_front = 1, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b1,     10'b1100_011100}, // D.28.3, disp_front = 1, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b0,     10'b0011_100010}, // D.29.3, disp_front = 1, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b0,     10'b0011_100001}, // D.30.3, disp_front = 1, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b0,     10'b0011_001010}, // D.31.3, disp_front = 1, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b1,     10'b1011_000110}, // D.00.4, disp_front = 1, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b1,     10'b1011_010001}, // D.01.4, disp_front = 1, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b1,     10'b1011_010010}, // D.02.4, disp_front = 1, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b0,     10'b0100_100011}, // D.03.4, disp_front = 1, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b1,     10'b1011_010100}, // D.04.4, disp_front = 1, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b0,     10'b0100_100101}, // D.05.4, disp_front = 1, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b0,     10'b0100_100110}, // D.06.4, disp_front = 1, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b0,     10'b0100_111000}, // D.07.4, disp_front = 1, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b1,     10'b1011_011000}, // D.08.4, disp_front = 1, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b0,     10'b0100_101001}, // D.09.4, disp_front = 1, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b0,     10'b0100_101010}, // D.10.4, disp_front = 1, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b0,     10'b0100_001011}, // D.11.4, disp_front = 1, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b0,     10'b0100_101100}, // D.12.4, disp_front = 1, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b0,     10'b0100_001101}, // D.13.4, disp_front = 1, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b0,     10'b0100_001110}, // D.14.4, disp_front = 1, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b1,     10'b1011_000101}, // D.15.4, disp_front = 1, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b1,     10'b1011_001001}, // D.16.4, disp_front = 1, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b0,     10'b0100_110001}, // D.17.4, disp_front = 1, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b0,     10'b0100_110010}, // D.18.4, disp_front = 1, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b0,     10'b0100_010011}, // D.19.4, disp_front = 1, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b0,     10'b0100_110100}, // D.20.4, disp_front = 1, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b0,     10'b0100_010101}, // D.21.4, disp_front = 1, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b0,     10'b0100_010110}, // D.22.4, disp_front = 1, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b1,     10'b1011_101000}, // D.23.4, disp_front = 1, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b1,     10'b1011_001100}, // D.24.4, disp_front = 1, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b0,     10'b0100_011001}, // D.25.4, disp_front = 1, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b0,     10'b0100_011010}, // D.26.4, disp_front = 1, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b1,     10'b1011_100100}, // D.27.4, disp_front = 1, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b0,     10'b0100_011100}, // D.28.4, disp_front = 1, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b1,     10'b1011_100010}, // D.29.4, disp_front = 1, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b1,     10'b1011_100001}, // D.30.4, disp_front = 1, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b1,     10'b1011_001010}, // D.31.4, disp_front = 1, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b0,     10'b0101_000110}, // D.00.5, disp_front = 1, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b0,     10'b0101_010001}, // D.01.5, disp_front = 1, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b0,     10'b0101_010010}, // D.02.5, disp_front = 1, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b1,     10'b0101_100011}, // D.03.5, disp_front = 1, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b0,     10'b0101_010100}, // D.04.5, disp_front = 1, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b1,     10'b0101_100101}, // D.05.5, disp_front = 1, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b1,     10'b0101_100110}, // D.06.5, disp_front = 1, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b1,     10'b0101_111000}, // D.07.5, disp_front = 1, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b0,     10'b0101_011000}, // D.08.5, disp_front = 1, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b1,     10'b0101_101001}, // D.09.5, disp_front = 1, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b1,     10'b0101_101010}, // D.10.5, disp_front = 1, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b1,     10'b0101_001011}, // D.11.5, disp_front = 1, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b1,     10'b0101_101100}, // D.12.5, disp_front = 1, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b1,     10'b0101_001101}, // D.13.5, disp_front = 1, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b1,     10'b0101_001110}, // D.14.5, disp_front = 1, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b0,     10'b0101_000101}, // D.15.5, disp_front = 1, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b0,     10'b0101_001001}, // D.16.5, disp_front = 1, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b1,     10'b0101_110001}, // D.17.5, disp_front = 1, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b1,     10'b0101_110010}, // D.18.5, disp_front = 1, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b1,     10'b0101_010011}, // D.19.5, disp_front = 1, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b1,     10'b0101_110100}, // D.20.5, disp_front = 1, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b1,     10'b0101_010101}, // D.21.5, disp_front = 1, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b1,     10'b0101_010110}, // D.22.5, disp_front = 1, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b0,     10'b0101_101000}, // D.23.5, disp_front = 1, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b0,     10'b0101_001100}, // D.24.5, disp_front = 1, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b1,     10'b0101_011001}, // D.25.5, disp_front = 1, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b1,     10'b0101_011010}, // D.26.5, disp_front = 1, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b0,     10'b0101_100100}, // D.27.5, disp_front = 1, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b1,     10'b0101_011100}, // D.28.5, disp_front = 1, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b0,     10'b0101_100010}, // D.29.5, disp_front = 1, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b0,     10'b0101_100001}, // D.30.5, disp_front = 1, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b0,     10'b0101_001010}, // D.31.5, disp_front = 1, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b0,     10'b0110_000110}, // D.00.6, disp_front = 1, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b0,     10'b0110_010001}, // D.01.6, disp_front = 1, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b0,     10'b0110_010010}, // D.02.6, disp_front = 1, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b1,     10'b0110_100011}, // D.03.6, disp_front = 1, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b0,     10'b0110_010100}, // D.04.6, disp_front = 1, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b1,     10'b0110_100101}, // D.05.6, disp_front = 1, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b1,     10'b0110_100110}, // D.06.6, disp_front = 1, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b1,     10'b0110_111000}, // D.07.6, disp_front = 1, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b0,     10'b0110_011000}, // D.08.6, disp_front = 1, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b1,     10'b0110_101001}, // D.09.6, disp_front = 1, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b1,     10'b0110_101010}, // D.10.6, disp_front = 1, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b1,     10'b0110_001011}, // D.11.6, disp_front = 1, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b1,     10'b0110_101100}, // D.12.6, disp_front = 1, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b1,     10'b0110_001101}, // D.13.6, disp_front = 1, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b1,     10'b0110_001110}, // D.14.6, disp_front = 1, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b0,     10'b0110_000101}, // D.15.6, disp_front = 1, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b0,     10'b0110_001001}, // D.16.6, disp_front = 1, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b1,     10'b0110_110001}, // D.17.6, disp_front = 1, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b1,     10'b0110_110010}, // D.18.6, disp_front = 1, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b1,     10'b0110_010011}, // D.19.6, disp_front = 1, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b1,     10'b0110_110100}, // D.20.6, disp_front = 1, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b1,     10'b0110_010101}, // D.21.6, disp_front = 1, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b1,     10'b0110_010110}, // D.22.6, disp_front = 1, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b0,     10'b0110_101000}, // D.23.6, disp_front = 1, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b0,     10'b0110_001100}, // D.24.6, disp_front = 1, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b1,     10'b0110_011001}, // D.25.6, disp_front = 1, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b1,     10'b0110_011010}, // D.26.6, disp_front = 1, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b0,     10'b0110_100100}, // D.27.6, disp_front = 1, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b1,     10'b0110_011100}, // D.28.6, disp_front = 1, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b0,     10'b0110_100010}, // D.29.6, disp_front = 1, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b0,     10'b0110_100001}, // D.30.6, disp_front = 1, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b0,     10'b0110_001010}, // D.31.6, disp_front = 1, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b1,     10'b0111_000110}, // D.00.7, disp_front = 1, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b1,     10'b0111_010001}, // D.01.7, disp_front = 1, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b1,     10'b0111_010010}, // D.02.7, disp_front = 1, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b0,     10'b1000_100011}, // D.03.7, disp_front = 1, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b1,     10'b0111_010100}, // D.04.7, disp_front = 1, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b0,     10'b1000_100101}, // D.05.7, disp_front = 1, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b0,     10'b1000_100110}, // D.06.7, disp_front = 1, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b0,     10'b1000_111000}, // D.07.7, disp_front = 1, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b1,     10'b0111_011000}, // D.08.7, disp_front = 1, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b0,     10'b1000_101001}, // D.09.7, disp_front = 1, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b0,     10'b1000_101010}, // D.10.7, disp_front = 1, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b0,     10'b0001_001011}, // D.11.7, disp_front = 1, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b0,     10'b1000_101100}, // D.12.7, disp_front = 1, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b0,     10'b0001_001101}, // D.13.7, disp_front = 1, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b0,     10'b0001_001110}, // D.14.7, disp_front = 1, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b1,     10'b0111_000101}, // D.15.7, disp_front = 1, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b1,     10'b0111_001001}, // D.16.7, disp_front = 1, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b0,     10'b1000_110001}, // D.17.7, disp_front = 1, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b0,     10'b1000_110010}, // D.18.7, disp_front = 1, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b0,     10'b1000_010011}, // D.19.7, disp_front = 1, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b0,     10'b1000_110100}, // D.20.7, disp_front = 1, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b0,     10'b1000_010101}, // D.21.7, disp_front = 1, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b0,     10'b1000_010110}, // D.22.7, disp_front = 1, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b1,     10'b0111_101000}, // D.23.7, disp_front = 1, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b1,     10'b0111_001100}, // D.24.7, disp_front = 1, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b0,     10'b1000_011001}, // D.25.7, disp_front = 1, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b0,     10'b1000_011010}, // D.26.7, disp_front = 1, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b1,     10'b0111_100100}, // D.27.7, disp_front = 1, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b0,     10'b1000_011100}, // D.28.7, disp_front = 1, K = 0 disp_end = 0, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b1,     10'b0111_100010}, // D.29.7, disp_front = 1, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b1,     10'b0111_100001}, // D.30.7, disp_front = 1, K = 0 disp_end = 1, code_err = 0
      {1'b0,      1'b1,       1'b0,     1'b1,     10'b0111_001010}, // D.31.7, disp_front = 1, K = 0 disp_end = 1, code_err = 0
      {1'b1,      1'b0,       1'b1,     1'b0,     10'b0010_111001}, // K.00.0, disp_front = 0, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b0,     10'b0010_101110}, // K.01.0, disp_front = 0, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b0,     10'b0010_101101}, // K.02.0, disp_front = 0, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b1,     10'b1101_100011}, // K.03.0, disp_front = 0, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b0,     10'b0010_101011}, // K.04.0, disp_front = 0, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b1,     10'b1101_100101}, // K.05.0, disp_front = 0, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b1,     10'b1101_100110}, // K.06.0, disp_front = 0, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b1,     10'b1101_000111}, // K.07.0, disp_front = 0, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b0,     10'b0010_100111}, // K.08.0, disp_front = 0, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b1,     10'b1101_101001}, // K.09.0, disp_front = 0, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b1,     10'b1101_101010}, // K.10.0, disp_front = 0, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b1,     10'b1101_001011}, // K.11.0, disp_front = 0, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b1,     10'b1101_101100}, // K.12.0, disp_front = 0, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b1,     10'b1101_001101}, // K.13.0, disp_front = 0, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b1,     10'b1101_001110}, // K.14.0, disp_front = 0, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b0,     10'b0010_111010}, // K.15.0, disp_front = 0, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b0,     10'b0010_110110}, // K.16.0, disp_front = 0, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b1,     10'b1101_110001}, // K.17.0, disp_front = 0, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b1,     10'b1101_110010}, // K.18.0, disp_front = 0, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b1,     10'b1101_010011}, // K.19.0, disp_front = 0, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b1,     10'b1101_110100}, // K.20.0, disp_front = 0, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b1,     10'b1101_010101}, // K.21.0, disp_front = 0, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b1,     10'b1101_010110}, // K.22.0, disp_front = 0, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b0,     10'b0010_010111}, // K.23.0, disp_front = 0, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b0,     10'b0010_110011}, // K.24.0, disp_front = 0, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b1,     10'b1101_011001}, // K.25.0, disp_front = 0, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b1,     10'b1101_011010}, // K.26.0, disp_front = 0, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b0,     10'b0010_011011}, // K.27.0, disp_front = 0, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b0,       1'b0,     1'b0,     10'b0010_111100}, // K.28.0, disp_front = 0, K = 1 disp_end = 0, code_err = 0
      {1'b1,      1'b0,       1'b1,     1'b0,     10'b0010_011101}, // K.29.0, disp_front = 0, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b0,     10'b0010_011110}, // K.30.0, disp_front = 0, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b0,     10'b0010_110101}, // K.31.0, disp_front = 0, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b1,     10'b1001_111001}, // K.00.1, disp_front = 0, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b1,     10'b1001_101110}, // K.01.1, disp_front = 0, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b1,     10'b1001_101101}, // K.02.1, disp_front = 0, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b0,     10'b0110_100011}, // K.03.1, disp_front = 0, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b1,     10'b1001_101011}, // K.04.1, disp_front = 0, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b0,     10'b0110_100101}, // K.05.1, disp_front = 0, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b0,     10'b0110_100110}, // K.06.1, disp_front = 0, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b0,     10'b0110_000111}, // K.07.1, disp_front = 0, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b1,     10'b1001_100111}, // K.08.1, disp_front = 0, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b0,     10'b0110_101001}, // K.09.1, disp_front = 0, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b0,     10'b0110_101010}, // K.10.1, disp_front = 0, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b0,     10'b0110_001011}, // K.11.1, disp_front = 0, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b0,     10'b0110_101100}, // K.12.1, disp_front = 0, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b0,     10'b0110_001101}, // K.13.1, disp_front = 0, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b0,     10'b0110_001110}, // K.14.1, disp_front = 0, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b1,     10'b1001_111010}, // K.15.1, disp_front = 0, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b1,     10'b1001_110110}, // K.16.1, disp_front = 0, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b0,     10'b0110_110001}, // K.17.1, disp_front = 0, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b0,     10'b0110_110010}, // K.18.1, disp_front = 0, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b0,     10'b0110_010011}, // K.19.1, disp_front = 0, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b0,     10'b0110_110100}, // K.20.1, disp_front = 0, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b0,     10'b0110_010101}, // K.21.1, disp_front = 0, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b0,     10'b0110_010110}, // K.22.1, disp_front = 0, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b1,     10'b1001_010111}, // K.23.1, disp_front = 0, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b1,     10'b1001_110011}, // K.24.1, disp_front = 0, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b0,     10'b0110_011001}, // K.25.1, disp_front = 0, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b0,     10'b0110_011010}, // K.26.1, disp_front = 0, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b1,     10'b1001_011011}, // K.27.1, disp_front = 0, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b0,       1'b0,     1'b1,     10'b1001_111100}, // K.28.1, disp_front = 0, K = 1 disp_end = 1, code_err = 0
      {1'b1,      1'b0,       1'b1,     1'b1,     10'b1001_011101}, // K.29.1, disp_front = 0, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b1,     10'b1001_011110}, // K.30.1, disp_front = 0, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b1,     10'b1001_110101}, // K.31.1, disp_front = 0, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b1,     10'b1010_111001}, // K.00.2, disp_front = 0, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b1,     10'b1010_101110}, // K.01.2, disp_front = 0, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b1,     10'b1010_101101}, // K.02.2, disp_front = 0, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b0,     10'b0101_100011}, // K.03.2, disp_front = 0, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b1,     10'b1010_101011}, // K.04.2, disp_front = 0, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b0,     10'b0101_100101}, // K.05.2, disp_front = 0, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b0,     10'b0101_100110}, // K.06.2, disp_front = 0, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b0,     10'b0101_000111}, // K.07.2, disp_front = 0, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b1,     10'b1010_100111}, // K.08.2, disp_front = 0, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b0,     10'b0101_101001}, // K.09.2, disp_front = 0, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b0,     10'b0101_101010}, // K.10.2, disp_front = 0, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b0,     10'b0101_001011}, // K.11.2, disp_front = 0, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b0,     10'b0101_101100}, // K.12.2, disp_front = 0, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b0,     10'b0101_001101}, // K.13.2, disp_front = 0, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b0,     10'b0101_001110}, // K.14.2, disp_front = 0, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b1,     10'b1010_111010}, // K.15.2, disp_front = 0, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b1,     10'b1010_110110}, // K.16.2, disp_front = 0, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b0,     10'b0101_110001}, // K.17.2, disp_front = 0, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b0,     10'b0101_110010}, // K.18.2, disp_front = 0, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b0,     10'b0101_010011}, // K.19.2, disp_front = 0, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b0,     10'b0101_110100}, // K.20.2, disp_front = 0, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b0,     10'b0101_010101}, // K.21.2, disp_front = 0, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b0,     10'b0101_010110}, // K.22.2, disp_front = 0, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b1,     10'b1010_010111}, // K.23.2, disp_front = 0, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b1,     10'b1010_110011}, // K.24.2, disp_front = 0, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b0,     10'b0101_011001}, // K.25.2, disp_front = 0, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b0,     10'b0101_011010}, // K.26.2, disp_front = 0, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b1,     10'b1010_011011}, // K.27.2, disp_front = 0, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b0,       1'b0,     1'b1,     10'b1010_111100}, // K.28.2, disp_front = 0, K = 1 disp_end = 1, code_err = 0
      {1'b1,      1'b0,       1'b1,     1'b1,     10'b1010_011101}, // K.29.2, disp_front = 0, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b1,     10'b1010_011110}, // K.30.2, disp_front = 0, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b1,     10'b1010_110101}, // K.31.2, disp_front = 0, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b1,     10'b1100_111001}, // K.00.3, disp_front = 0, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b1,     10'b1100_101110}, // K.01.3, disp_front = 0, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b1,     10'b1100_101101}, // K.02.3, disp_front = 0, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b0,     10'b0011_100011}, // K.03.3, disp_front = 0, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b1,     10'b1100_101011}, // K.04.3, disp_front = 0, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b0,     10'b0011_100101}, // K.05.3, disp_front = 0, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b0,     10'b0011_100110}, // K.06.3, disp_front = 0, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b0,     10'b0011_000111}, // K.07.3, disp_front = 0, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b1,     10'b1100_100111}, // K.08.3, disp_front = 0, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b0,     10'b0011_101001}, // K.09.3, disp_front = 0, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b0,     10'b0011_101010}, // K.10.3, disp_front = 0, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b0,     10'b0011_001011}, // K.11.3, disp_front = 0, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b0,     10'b0011_101100}, // K.12.3, disp_front = 0, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b0,     10'b0011_001101}, // K.13.3, disp_front = 0, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b0,     10'b0011_001110}, // K.14.3, disp_front = 0, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b1,     10'b1100_111010}, // K.15.3, disp_front = 0, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b1,     10'b1100_110110}, // K.16.3, disp_front = 0, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b0,     10'b0011_110001}, // K.17.3, disp_front = 0, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b0,     10'b0011_110010}, // K.18.3, disp_front = 0, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b0,     10'b0011_010011}, // K.19.3, disp_front = 0, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b0,     10'b0011_110100}, // K.20.3, disp_front = 0, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b0,     10'b0011_010101}, // K.21.3, disp_front = 0, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b0,     10'b0011_010110}, // K.22.3, disp_front = 0, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b1,     10'b1100_010111}, // K.23.3, disp_front = 0, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b1,     10'b1100_110011}, // K.24.3, disp_front = 0, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b0,     10'b0011_011001}, // K.25.3, disp_front = 0, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b0,     10'b0011_011010}, // K.26.3, disp_front = 0, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b1,     10'b1100_011011}, // K.27.3, disp_front = 0, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b0,       1'b0,     1'b1,     10'b1100_111100}, // K.28.3, disp_front = 0, K = 1 disp_end = 1, code_err = 0
      {1'b1,      1'b0,       1'b1,     1'b1,     10'b1100_011101}, // K.29.3, disp_front = 0, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b1,     10'b1100_011110}, // K.30.3, disp_front = 0, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b1,     10'b1100_110101}, // K.31.3, disp_front = 0, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b0,     10'b0100_111001}, // K.00.4, disp_front = 0, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b0,     10'b0100_101110}, // K.01.4, disp_front = 0, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b0,     10'b0100_101101}, // K.02.4, disp_front = 0, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b1,     10'b1011_100011}, // K.03.4, disp_front = 0, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b0,     10'b0100_101011}, // K.04.4, disp_front = 0, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b1,     10'b1011_100101}, // K.05.4, disp_front = 0, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b1,     10'b1011_100110}, // K.06.4, disp_front = 0, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b1,     10'b1011_000111}, // K.07.4, disp_front = 0, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b0,     10'b0100_100111}, // K.08.4, disp_front = 0, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b1,     10'b1011_101001}, // K.09.4, disp_front = 0, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b1,     10'b1011_101010}, // K.10.4, disp_front = 0, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b1,     10'b1011_001011}, // K.11.4, disp_front = 0, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b1,     10'b1011_101100}, // K.12.4, disp_front = 0, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b1,     10'b1011_001101}, // K.13.4, disp_front = 0, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b1,     10'b1011_001110}, // K.14.4, disp_front = 0, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b0,     10'b0100_111010}, // K.15.4, disp_front = 0, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b0,     10'b0100_110110}, // K.16.4, disp_front = 0, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b1,     10'b1011_110001}, // K.17.4, disp_front = 0, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b1,     10'b1011_110010}, // K.18.4, disp_front = 0, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b1,     10'b1011_010011}, // K.19.4, disp_front = 0, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b1,     10'b1011_110100}, // K.20.4, disp_front = 0, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b1,     10'b1011_010101}, // K.21.4, disp_front = 0, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b1,     10'b1011_010110}, // K.22.4, disp_front = 0, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b0,     10'b0100_010111}, // K.23.4, disp_front = 0, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b0,     10'b0100_110011}, // K.24.4, disp_front = 0, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b1,     10'b1011_011001}, // K.25.4, disp_front = 0, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b1,     10'b1011_011010}, // K.26.4, disp_front = 0, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b0,     10'b0100_011011}, // K.27.4, disp_front = 0, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b0,       1'b0,     1'b0,     10'b0100_111100}, // K.28.4, disp_front = 0, K = 1 disp_end = 0, code_err = 0
      {1'b1,      1'b0,       1'b1,     1'b0,     10'b0100_011101}, // K.29.4, disp_front = 0, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b0,     10'b0100_011110}, // K.30.4, disp_front = 0, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b0,     10'b0100_110101}, // K.31.4, disp_front = 0, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b1,     10'b0101_111001}, // K.00.5, disp_front = 0, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b1,     10'b0101_101110}, // K.01.5, disp_front = 0, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b1,     10'b0101_101101}, // K.02.5, disp_front = 0, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b0,     10'b1010_100011}, // K.03.5, disp_front = 0, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b1,     10'b0101_101011}, // K.04.5, disp_front = 0, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b0,     10'b1010_100101}, // K.05.5, disp_front = 0, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b0,     10'b1010_100110}, // K.06.5, disp_front = 0, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b0,     10'b1010_000111}, // K.07.5, disp_front = 0, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b1,     10'b0101_100111}, // K.08.5, disp_front = 0, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b0,     10'b1010_101001}, // K.09.5, disp_front = 0, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b0,     10'b1010_101010}, // K.10.5, disp_front = 0, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b0,     10'b1010_001011}, // K.11.5, disp_front = 0, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b0,     10'b1010_101100}, // K.12.5, disp_front = 0, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b0,     10'b1010_001101}, // K.13.5, disp_front = 0, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b0,     10'b1010_001110}, // K.14.5, disp_front = 0, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b1,     10'b0101_111010}, // K.15.5, disp_front = 0, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b1,     10'b0101_110110}, // K.16.5, disp_front = 0, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b0,     10'b1010_110001}, // K.17.5, disp_front = 0, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b0,     10'b1010_110010}, // K.18.5, disp_front = 0, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b0,     10'b1010_010011}, // K.19.5, disp_front = 0, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b0,     10'b1010_110100}, // K.20.5, disp_front = 0, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b0,     10'b1010_010101}, // K.21.5, disp_front = 0, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b0,     10'b1010_010110}, // K.22.5, disp_front = 0, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b1,     10'b0101_010111}, // K.23.5, disp_front = 0, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b1,     10'b0101_110011}, // K.24.5, disp_front = 0, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b0,     10'b1010_011001}, // K.25.5, disp_front = 0, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b0,     10'b1010_011010}, // K.26.5, disp_front = 0, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b1,     10'b0101_011011}, // K.27.5, disp_front = 0, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b0,       1'b0,     1'b1,     10'b0101_111100}, // K.28.5, disp_front = 0, K = 1 disp_end = 1, code_err = 0
      {1'b1,      1'b0,       1'b1,     1'b1,     10'b0101_011101}, // K.29.5, disp_front = 0, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b1,     10'b0101_011110}, // K.30.5, disp_front = 0, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b1,     10'b0101_110101}, // K.31.5, disp_front = 0, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b1,     10'b0110_111001}, // K.00.6, disp_front = 0, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b1,     10'b0110_101110}, // K.01.6, disp_front = 0, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b1,     10'b0110_101101}, // K.02.6, disp_front = 0, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b0,     10'b1001_100011}, // K.03.6, disp_front = 0, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b1,     10'b0110_101011}, // K.04.6, disp_front = 0, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b0,     10'b1001_100101}, // K.05.6, disp_front = 0, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b0,     10'b1001_100110}, // K.06.6, disp_front = 0, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b0,     10'b1001_000111}, // K.07.6, disp_front = 0, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b1,     10'b0110_100111}, // K.08.6, disp_front = 0, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b0,     10'b1001_101001}, // K.09.6, disp_front = 0, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b0,     10'b1001_101010}, // K.10.6, disp_front = 0, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b0,     10'b1001_001011}, // K.11.6, disp_front = 0, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b0,     10'b1001_101100}, // K.12.6, disp_front = 0, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b0,     10'b1001_001101}, // K.13.6, disp_front = 0, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b0,     10'b1001_001110}, // K.14.6, disp_front = 0, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b1,     10'b0110_111010}, // K.15.6, disp_front = 0, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b1,     10'b0110_110110}, // K.16.6, disp_front = 0, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b0,     10'b1001_110001}, // K.17.6, disp_front = 0, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b0,     10'b1001_110010}, // K.18.6, disp_front = 0, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b0,     10'b1001_010011}, // K.19.6, disp_front = 0, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b0,     10'b1001_110100}, // K.20.6, disp_front = 0, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b0,     10'b1001_010101}, // K.21.6, disp_front = 0, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b0,     10'b1001_010110}, // K.22.6, disp_front = 0, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b1,     10'b0110_010111}, // K.23.6, disp_front = 0, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b1,     10'b0110_110011}, // K.24.6, disp_front = 0, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b0,     10'b1001_011001}, // K.25.6, disp_front = 0, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b0,     10'b1001_011010}, // K.26.6, disp_front = 0, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b1,     10'b0110_011011}, // K.27.6, disp_front = 0, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b0,       1'b0,     1'b1,     10'b0110_111100}, // K.28.6, disp_front = 0, K = 1 disp_end = 1, code_err = 0
      {1'b1,      1'b0,       1'b1,     1'b1,     10'b0110_011101}, // K.29.6, disp_front = 0, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b1,     10'b0110_011110}, // K.30.6, disp_front = 0, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b1,     10'b0110_110101}, // K.31.6, disp_front = 0, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b0,     10'b0001_111001}, // K.00.7, disp_front = 0, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b0,     10'b0001_101110}, // K.01.7, disp_front = 0, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b0,     10'b0001_101101}, // K.02.7, disp_front = 0, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b1,     10'b1110_100011}, // K.03.7, disp_front = 0, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b0,     10'b0001_101011}, // K.04.7, disp_front = 0, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b1,     10'b1110_100101}, // K.05.7, disp_front = 0, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b1,     10'b1110_100110}, // K.06.7, disp_front = 0, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b1,     10'b1110_000111}, // K.07.7, disp_front = 0, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b0,     10'b0001_100111}, // K.08.7, disp_front = 0, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b1,     10'b1110_101001}, // K.09.7, disp_front = 0, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b1,     10'b1110_101010}, // K.10.7, disp_front = 0, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b1,     10'b1110_001011}, // K.11.7, disp_front = 0, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b1,     10'b1110_101100}, // K.12.7, disp_front = 0, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b1,     10'b1110_001101}, // K.13.7, disp_front = 0, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b1,     10'b1110_001110}, // K.14.7, disp_front = 0, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b0,     10'b0001_111010}, // K.15.7, disp_front = 0, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b0,     10'b0001_110110}, // K.16.7, disp_front = 0, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b1,     10'b1110_110001}, // K.17.7, disp_front = 0, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b1,     10'b1110_110010}, // K.18.7, disp_front = 0, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b1,     10'b1110_010011}, // K.19.7, disp_front = 0, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b1,     10'b1110_110100}, // K.20.7, disp_front = 0, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b1,     10'b1110_010101}, // K.21.7, disp_front = 0, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b1,     10'b1110_010110}, // K.22.7, disp_front = 0, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b0,       1'b0,     1'b0,     10'b0001_010111}, // K.23.7, disp_front = 0, K = 1 disp_end = 0, code_err = 0
      {1'b1,      1'b0,       1'b1,     1'b0,     10'b0001_110011}, // K.24.7, disp_front = 0, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b1,     10'b1110_011001}, // K.25.7, disp_front = 0, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b0,       1'b1,     1'b1,     10'b1110_011010}, // K.26.7, disp_front = 0, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b0,       1'b0,     1'b0,     10'b0001_011011}, // K.27.7, disp_front = 0, K = 1 disp_end = 0, code_err = 0
      {1'b1,      1'b0,       1'b0,     1'b0,     10'b0001_111100}, // K.28.7, disp_front = 0, K = 1 disp_end = 0, code_err = 0
      {1'b1,      1'b0,       1'b0,     1'b0,     10'b0001_011101}, // K.29.7, disp_front = 0, K = 1 disp_end = 0, code_err = 0
      {1'b1,      1'b0,       1'b0,     1'b0,     10'b0001_011110}, // K.30.7, disp_front = 0, K = 1 disp_end = 0, code_err = 0
      {1'b1,      1'b0,       1'b1,     1'b0,     10'b0001_110101}, // K.31.7, disp_front = 0, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b1,     10'b1101_000110}, // K.00.0, disp_front = 1, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b1,     10'b1101_010001}, // K.01.0, disp_front = 1, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b1,     10'b1101_010010}, // K.02.0, disp_front = 1, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b0,     10'b0010_100011}, // K.03.0, disp_front = 1, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b1,     10'b1101_010100}, // K.04.0, disp_front = 1, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b0,     10'b0010_100101}, // K.05.0, disp_front = 1, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b0,     10'b0010_100110}, // K.06.0, disp_front = 1, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b0,     10'b0010_111000}, // K.07.0, disp_front = 1, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b1,     10'b1101_011000}, // K.08.0, disp_front = 1, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b0,     10'b0010_101001}, // K.09.0, disp_front = 1, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b0,     10'b0010_101010}, // K.10.0, disp_front = 1, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b0,     10'b0010_001011}, // K.11.0, disp_front = 1, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b0,     10'b0010_101100}, // K.12.0, disp_front = 1, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b0,     10'b0010_001101}, // K.13.0, disp_front = 1, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b0,     10'b0010_001110}, // K.14.0, disp_front = 1, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b1,     10'b1101_000101}, // K.15.0, disp_front = 1, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b1,     10'b1101_001001}, // K.16.0, disp_front = 1, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b0,     10'b0010_110001}, // K.17.0, disp_front = 1, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b0,     10'b0010_110010}, // K.18.0, disp_front = 1, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b0,     10'b0010_010011}, // K.19.0, disp_front = 1, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b0,     10'b0010_110100}, // K.20.0, disp_front = 1, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b0,     10'b0010_010101}, // K.21.0, disp_front = 1, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b0,     10'b0010_010110}, // K.22.0, disp_front = 1, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b1,     10'b1101_101000}, // K.23.0, disp_front = 1, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b1,     10'b1101_001100}, // K.24.0, disp_front = 1, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b0,     10'b0010_011001}, // K.25.0, disp_front = 1, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b0,     10'b0010_011010}, // K.26.0, disp_front = 1, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b1,     10'b1101_100100}, // K.27.0, disp_front = 1, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b1,       1'b0,     1'b1,     10'b1101_000011}, // K.28.0, disp_front = 1, K = 1 disp_end = 1, code_err = 0
      {1'b1,      1'b1,       1'b1,     1'b1,     10'b1101_100010}, // K.29.0, disp_front = 1, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b1,     10'b1101_100001}, // K.30.0, disp_front = 1, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b1,     10'b1101_001010}, // K.31.0, disp_front = 1, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b0,     10'b0110_000110}, // K.00.1, disp_front = 1, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b0,     10'b0110_010001}, // K.01.1, disp_front = 1, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b0,     10'b0110_010010}, // K.02.1, disp_front = 1, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b1,     10'b1001_100011}, // K.03.1, disp_front = 1, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b0,     10'b0110_010100}, // K.04.1, disp_front = 1, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b1,     10'b1001_100101}, // K.05.1, disp_front = 1, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b1,     10'b1001_100110}, // K.06.1, disp_front = 1, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b1,     10'b1001_111000}, // K.07.1, disp_front = 1, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b0,     10'b0110_011000}, // K.08.1, disp_front = 1, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b1,     10'b1001_101001}, // K.09.1, disp_front = 1, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b1,     10'b1001_101010}, // K.10.1, disp_front = 1, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b1,     10'b1001_001011}, // K.11.1, disp_front = 1, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b1,     10'b1001_101100}, // K.12.1, disp_front = 1, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b1,     10'b1001_001101}, // K.13.1, disp_front = 1, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b1,     10'b1001_001110}, // K.14.1, disp_front = 1, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b0,     10'b0110_000101}, // K.15.1, disp_front = 1, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b0,     10'b0110_001001}, // K.16.1, disp_front = 1, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b1,     10'b1001_110001}, // K.17.1, disp_front = 1, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b1,     10'b1001_110010}, // K.18.1, disp_front = 1, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b1,     10'b1001_010011}, // K.19.1, disp_front = 1, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b1,     10'b1001_110100}, // K.20.1, disp_front = 1, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b1,     10'b1001_010101}, // K.21.1, disp_front = 1, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b1,     10'b1001_010110}, // K.22.1, disp_front = 1, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b0,     10'b0110_101000}, // K.23.1, disp_front = 1, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b0,     10'b0110_001100}, // K.24.1, disp_front = 1, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b1,     10'b1001_011001}, // K.25.1, disp_front = 1, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b1,     10'b1001_011010}, // K.26.1, disp_front = 1, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b0,     10'b0110_100100}, // K.27.1, disp_front = 1, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b1,       1'b0,     1'b0,     10'b0110_000011}, // K.28.1, disp_front = 1, K = 1 disp_end = 0, code_err = 0
      {1'b1,      1'b1,       1'b1,     1'b0,     10'b0110_100010}, // K.29.1, disp_front = 1, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b0,     10'b0110_100001}, // K.30.1, disp_front = 1, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b0,     10'b0110_001010}, // K.31.1, disp_front = 1, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b0,     10'b0101_000110}, // K.00.2, disp_front = 1, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b0,     10'b0101_010001}, // K.01.2, disp_front = 1, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b0,     10'b0101_010010}, // K.02.2, disp_front = 1, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b1,     10'b1010_100011}, // K.03.2, disp_front = 1, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b0,     10'b0101_010100}, // K.04.2, disp_front = 1, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b1,     10'b1010_100101}, // K.05.2, disp_front = 1, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b1,     10'b1010_100110}, // K.06.2, disp_front = 1, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b1,     10'b1010_111000}, // K.07.2, disp_front = 1, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b0,     10'b0101_011000}, // K.08.2, disp_front = 1, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b1,     10'b1010_101001}, // K.09.2, disp_front = 1, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b1,     10'b1010_101010}, // K.10.2, disp_front = 1, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b1,     10'b1010_001011}, // K.11.2, disp_front = 1, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b1,     10'b1010_101100}, // K.12.2, disp_front = 1, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b1,     10'b1010_001101}, // K.13.2, disp_front = 1, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b1,     10'b1010_001110}, // K.14.2, disp_front = 1, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b0,     10'b0101_000101}, // K.15.2, disp_front = 1, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b0,     10'b0101_001001}, // K.16.2, disp_front = 1, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b1,     10'b1010_110001}, // K.17.2, disp_front = 1, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b1,     10'b1010_110010}, // K.18.2, disp_front = 1, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b1,     10'b1010_010011}, // K.19.2, disp_front = 1, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b1,     10'b1010_110100}, // K.20.2, disp_front = 1, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b1,     10'b1010_010101}, // K.21.2, disp_front = 1, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b1,     10'b1010_010110}, // K.22.2, disp_front = 1, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b0,     10'b0101_101000}, // K.23.2, disp_front = 1, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b0,     10'b0101_001100}, // K.24.2, disp_front = 1, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b1,     10'b1010_011001}, // K.25.2, disp_front = 1, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b1,     10'b1010_011010}, // K.26.2, disp_front = 1, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b0,     10'b0101_100100}, // K.27.2, disp_front = 1, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b1,       1'b0,     1'b0,     10'b0101_000011}, // K.28.2, disp_front = 1, K = 1 disp_end = 0, code_err = 0
      {1'b1,      1'b1,       1'b1,     1'b0,     10'b0101_100010}, // K.29.2, disp_front = 1, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b0,     10'b0101_100001}, // K.30.2, disp_front = 1, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b0,     10'b0101_001010}, // K.31.2, disp_front = 1, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b0,     10'b0011_000110}, // K.00.3, disp_front = 1, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b0,     10'b0011_010001}, // K.01.3, disp_front = 1, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b0,     10'b0011_010010}, // K.02.3, disp_front = 1, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b1,     10'b1100_100011}, // K.03.3, disp_front = 1, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b0,     10'b0011_010100}, // K.04.3, disp_front = 1, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b1,     10'b1100_100101}, // K.05.3, disp_front = 1, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b1,     10'b1100_100110}, // K.06.3, disp_front = 1, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b1,     10'b1100_111000}, // K.07.3, disp_front = 1, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b0,     10'b0011_011000}, // K.08.3, disp_front = 1, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b1,     10'b1100_101001}, // K.09.3, disp_front = 1, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b1,     10'b1100_101010}, // K.10.3, disp_front = 1, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b1,     10'b1100_001011}, // K.11.3, disp_front = 1, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b1,     10'b1100_101100}, // K.12.3, disp_front = 1, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b1,     10'b1100_001101}, // K.13.3, disp_front = 1, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b1,     10'b1100_001110}, // K.14.3, disp_front = 1, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b0,     10'b0011_000101}, // K.15.3, disp_front = 1, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b0,     10'b0011_001001}, // K.16.3, disp_front = 1, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b1,     10'b1100_110001}, // K.17.3, disp_front = 1, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b1,     10'b1100_110010}, // K.18.3, disp_front = 1, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b1,     10'b1100_010011}, // K.19.3, disp_front = 1, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b1,     10'b1100_110100}, // K.20.3, disp_front = 1, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b1,     10'b1100_010101}, // K.21.3, disp_front = 1, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b1,     10'b1100_010110}, // K.22.3, disp_front = 1, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b0,     10'b0011_101000}, // K.23.3, disp_front = 1, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b0,     10'b0011_001100}, // K.24.3, disp_front = 1, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b1,     10'b1100_011001}, // K.25.3, disp_front = 1, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b1,     10'b1100_011010}, // K.26.3, disp_front = 1, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b0,     10'b0011_100100}, // K.27.3, disp_front = 1, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b1,       1'b0,     1'b0,     10'b0011_000011}, // K.28.3, disp_front = 1, K = 1 disp_end = 0, code_err = 0
      {1'b1,      1'b1,       1'b1,     1'b0,     10'b0011_100010}, // K.29.3, disp_front = 1, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b0,     10'b0011_100001}, // K.30.3, disp_front = 1, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b0,     10'b0011_001010}, // K.31.3, disp_front = 1, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b1,     10'b1011_000110}, // K.00.4, disp_front = 1, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b1,     10'b1011_010001}, // K.01.4, disp_front = 1, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b1,     10'b1011_010010}, // K.02.4, disp_front = 1, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b0,     10'b0100_100011}, // K.03.4, disp_front = 1, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b1,     10'b1011_010100}, // K.04.4, disp_front = 1, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b0,     10'b0100_100101}, // K.05.4, disp_front = 1, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b0,     10'b0100_100110}, // K.06.4, disp_front = 1, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b0,     10'b0100_111000}, // K.07.4, disp_front = 1, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b1,     10'b1011_011000}, // K.08.4, disp_front = 1, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b0,     10'b0100_101001}, // K.09.4, disp_front = 1, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b0,     10'b0100_101010}, // K.10.4, disp_front = 1, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b0,     10'b0100_001011}, // K.11.4, disp_front = 1, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b0,     10'b0100_101100}, // K.12.4, disp_front = 1, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b0,     10'b0100_001101}, // K.13.4, disp_front = 1, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b0,     10'b0100_001110}, // K.14.4, disp_front = 1, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b1,     10'b1011_000101}, // K.15.4, disp_front = 1, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b1,     10'b1011_001001}, // K.16.4, disp_front = 1, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b0,     10'b0100_110001}, // K.17.4, disp_front = 1, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b0,     10'b0100_110010}, // K.18.4, disp_front = 1, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b0,     10'b0100_010011}, // K.19.4, disp_front = 1, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b0,     10'b0100_110100}, // K.20.4, disp_front = 1, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b0,     10'b0100_010101}, // K.21.4, disp_front = 1, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b0,     10'b0100_010110}, // K.22.4, disp_front = 1, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b1,     10'b1011_101000}, // K.23.4, disp_front = 1, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b1,     10'b1011_001100}, // K.24.4, disp_front = 1, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b0,     10'b0100_011001}, // K.25.4, disp_front = 1, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b0,     10'b0100_011010}, // K.26.4, disp_front = 1, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b1,     10'b1011_100100}, // K.27.4, disp_front = 1, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b1,       1'b0,     1'b1,     10'b1011_000011}, // K.28.4, disp_front = 1, K = 1 disp_end = 1, code_err = 0
      {1'b1,      1'b1,       1'b1,     1'b1,     10'b1011_100010}, // K.29.4, disp_front = 1, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b1,     10'b1011_100001}, // K.30.4, disp_front = 1, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b1,     10'b1011_001010}, // K.31.4, disp_front = 1, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b0,     10'b1010_000110}, // K.00.5, disp_front = 1, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b0,     10'b1010_010001}, // K.01.5, disp_front = 1, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b0,     10'b1010_010010}, // K.02.5, disp_front = 1, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b1,     10'b0101_100011}, // K.03.5, disp_front = 1, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b0,     10'b1010_010100}, // K.04.5, disp_front = 1, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b1,     10'b0101_100101}, // K.05.5, disp_front = 1, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b1,     10'b0101_100110}, // K.06.5, disp_front = 1, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b1,     10'b0101_111000}, // K.07.5, disp_front = 1, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b0,     10'b1010_011000}, // K.08.5, disp_front = 1, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b1,     10'b0101_101001}, // K.09.5, disp_front = 1, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b1,     10'b0101_101010}, // K.10.5, disp_front = 1, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b1,     10'b0101_001011}, // K.11.5, disp_front = 1, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b1,     10'b0101_101100}, // K.12.5, disp_front = 1, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b1,     10'b0101_001101}, // K.13.5, disp_front = 1, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b1,     10'b0101_001110}, // K.14.5, disp_front = 1, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b0,     10'b1010_000101}, // K.15.5, disp_front = 1, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b0,     10'b1010_001001}, // K.16.5, disp_front = 1, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b1,     10'b0101_110001}, // K.17.5, disp_front = 1, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b1,     10'b0101_110010}, // K.18.5, disp_front = 1, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b1,     10'b0101_010011}, // K.19.5, disp_front = 1, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b1,     10'b0101_110100}, // K.20.5, disp_front = 1, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b1,     10'b0101_010101}, // K.21.5, disp_front = 1, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b1,     10'b0101_010110}, // K.22.5, disp_front = 1, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b0,     10'b1010_101000}, // K.23.5, disp_front = 1, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b0,     10'b1010_001100}, // K.24.5, disp_front = 1, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b1,     10'b0101_011001}, // K.25.5, disp_front = 1, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b1,     10'b0101_011010}, // K.26.5, disp_front = 1, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b0,     10'b1010_100100}, // K.27.5, disp_front = 1, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b1,       1'b0,     1'b0,     10'b1010_000011}, // K.28.5, disp_front = 1, K = 1 disp_end = 0, code_err = 0
      {1'b1,      1'b1,       1'b1,     1'b0,     10'b1010_100010}, // K.29.5, disp_front = 1, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b0,     10'b1010_100001}, // K.30.5, disp_front = 1, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b0,     10'b1010_001010}, // K.31.5, disp_front = 1, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b0,     10'b1001_000110}, // K.00.6, disp_front = 1, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b0,     10'b1001_010001}, // K.01.6, disp_front = 1, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b0,     10'b1001_010010}, // K.02.6, disp_front = 1, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b1,     10'b0110_100011}, // K.03.6, disp_front = 1, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b0,     10'b1001_010100}, // K.04.6, disp_front = 1, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b1,     10'b0110_100101}, // K.05.6, disp_front = 1, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b1,     10'b0110_100110}, // K.06.6, disp_front = 1, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b1,     10'b0110_111000}, // K.07.6, disp_front = 1, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b0,     10'b1001_011000}, // K.08.6, disp_front = 1, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b1,     10'b0110_101001}, // K.09.6, disp_front = 1, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b1,     10'b0110_101010}, // K.10.6, disp_front = 1, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b1,     10'b0110_001011}, // K.11.6, disp_front = 1, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b1,     10'b0110_101100}, // K.12.6, disp_front = 1, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b1,     10'b0110_001101}, // K.13.6, disp_front = 1, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b1,     10'b0110_001110}, // K.14.6, disp_front = 1, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b0,     10'b1001_000101}, // K.15.6, disp_front = 1, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b0,     10'b1001_001001}, // K.16.6, disp_front = 1, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b1,     10'b0110_110001}, // K.17.6, disp_front = 1, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b1,     10'b0110_110010}, // K.18.6, disp_front = 1, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b1,     10'b0110_010011}, // K.19.6, disp_front = 1, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b1,     10'b0110_110100}, // K.20.6, disp_front = 1, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b1,     10'b0110_010101}, // K.21.6, disp_front = 1, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b1,     10'b0110_010110}, // K.22.6, disp_front = 1, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b0,     10'b1001_101000}, // K.23.6, disp_front = 1, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b0,     10'b1001_001100}, // K.24.6, disp_front = 1, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b1,     10'b0110_011001}, // K.25.6, disp_front = 1, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b1,     10'b0110_011010}, // K.26.6, disp_front = 1, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b0,     10'b1001_100100}, // K.27.6, disp_front = 1, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b1,       1'b0,     1'b0,     10'b1001_000011}, // K.28.6, disp_front = 1, K = 1 disp_end = 0, code_err = 0
      {1'b1,      1'b1,       1'b1,     1'b0,     10'b1001_100010}, // K.29.6, disp_front = 1, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b0,     10'b1001_100001}, // K.30.6, disp_front = 1, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b0,     10'b1001_001010}, // K.31.6, disp_front = 1, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b1,     10'b1110_000110}, // K.00.7, disp_front = 1, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b1,     10'b1110_010001}, // K.01.7, disp_front = 1, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b1,     10'b1110_010010}, // K.02.7, disp_front = 1, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b0,     10'b0001_100011}, // K.03.7, disp_front = 1, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b1,     10'b1110_010100}, // K.04.7, disp_front = 1, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b0,     10'b0001_100101}, // K.05.7, disp_front = 1, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b0,     10'b0001_100110}, // K.06.7, disp_front = 1, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b0,     10'b0001_111000}, // K.07.7, disp_front = 1, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b1,     10'b1110_011000}, // K.08.7, disp_front = 1, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b0,     10'b0001_101001}, // K.09.7, disp_front = 1, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b0,     10'b0001_101010}, // K.10.7, disp_front = 1, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b0,     10'b0001_001011}, // K.11.7, disp_front = 1, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b0,     10'b0001_101100}, // K.12.7, disp_front = 1, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b0,     10'b0001_001101}, // K.13.7, disp_front = 1, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b0,     10'b0001_001110}, // K.14.7, disp_front = 1, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b1,     10'b1110_000101}, // K.15.7, disp_front = 1, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b1,     10'b1110_001001}, // K.16.7, disp_front = 1, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b0,     10'b0001_110001}, // K.17.7, disp_front = 1, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b0,     10'b0001_110010}, // K.18.7, disp_front = 1, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b0,     10'b0001_010011}, // K.19.7, disp_front = 1, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b0,     10'b0001_110100}, // K.20.7, disp_front = 1, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b0,     10'b0001_010101}, // K.21.7, disp_front = 1, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b0,     10'b0001_010110}, // K.22.7, disp_front = 1, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b1,       1'b0,     1'b1,     10'b1110_101000}, // K.23.7, disp_front = 1, K = 1 disp_end = 1, code_err = 0
      {1'b1,      1'b1,       1'b1,     1'b1,     10'b1110_001100}, // K.24.7, disp_front = 1, K = 1 disp_end = 1, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b0,     10'b0001_011001}, // K.25.7, disp_front = 1, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b1,       1'b1,     1'b0,     10'b0001_011010}, // K.26.7, disp_front = 1, K = 1 disp_end = 0, code_err = 1
      {1'b1,      1'b1,       1'b0,     1'b1,     10'b1110_100100}, // K.27.7, disp_front = 1, K = 1 disp_end = 1, code_err = 0
      {1'b1,      1'b1,       1'b0,     1'b1,     10'b1110_000011}, // K.28.7, disp_front = 1, K = 1 disp_end = 1, code_err = 0
      {1'b1,      1'b1,       1'b0,     1'b1,     10'b1110_100010}, // K.29.7, disp_front = 1, K = 1 disp_end = 1, code_err = 0
      {1'b1,      1'b1,       1'b0,     1'b1,     10'b1110_100001}, // K.30.7, disp_front = 1, K = 1 disp_end = 1, code_err = 0
      {1'b1,      1'b1,       1'b1,     1'b1,     10'b1110_001010}  // K.31.7, disp_front = 1, K = 1 disp_end = 1, code_err = 1
  };

endpackage