package dec_10b8b_pkg;

  logic [12:0] dec_symb [0:2047] = '{
    //disp_front  disp_err  code_err  ctrl_symb disp_end  octet
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b0,     8'b00000000}, // D.00.0, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b0,     8'b00000000}, // D.00.0, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b0,     8'b00000000}, // D.00.0, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b0,     8'b00011100}, // D.28.0, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b0,     8'b00000000}, // D.00.0, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b0,     8'b00001111}, // D.15.0, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b0,     8'b00000000}, // D.00.0, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b1,     8'b00000111}, // D.07.0, disp_front = 0, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b0,     8'b00000000}, // D.00.0, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b0,     8'b00010000}, // D.16.0, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b0,     8'b00011111}, // D.31.0, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b1,     8'b00001011}, // D.11.0, disp_front = 0, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b0,     8'b00011000}, // D.24.0, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b1,     8'b00001101}, // D.13.0, disp_front = 0, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b1,     8'b00001110}, // D.14.0, disp_front = 0, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b0,     8'b00000000}, // D.00.0, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b0,     8'b00000000}, // D.00.0, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b0,     8'b00000001}, // D.01.0, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b0,     8'b00000010}, // D.02.0, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b1,     8'b00010011}, // D.19.0, disp_front = 0, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b0,     8'b00000100}, // D.04.0, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b1,     8'b00010101}, // D.21.0, disp_front = 0, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b1,     8'b00010110}, // D.22.0, disp_front = 0, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b0,     8'b00010111}, // D.23.0, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b0,     8'b00001000}, // D.08.0, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b1,     8'b00011001}, // D.25.0, disp_front = 0, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b1,     8'b00011010}, // D.26.0, disp_front = 0, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b0,     8'b00011011}, // D.27.0, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b1,     8'b00011100}, // D.28.0, disp_front = 0, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b0,     8'b00011101}, // D.29.0, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b0,     8'b00011110}, // D.30.0, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b0,     8'b00000000}, // D.00.0, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b0,     8'b00000000}, // D.00.0, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b0,     8'b00011110}, // D.30.0, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b0,     8'b00011101}, // D.29.0, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b1,     8'b00000011}, // D.03.0, disp_front = 0, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b0,     8'b00011011}, // D.27.0, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b1,     8'b00000101}, // D.05.0, disp_front = 0, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b1,     8'b00000110}, // D.06.0, disp_front = 0, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b0,     8'b00001000}, // D.08.0, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b0,     8'b00010111}, // D.23.0, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b1,     8'b00001001}, // D.09.0, disp_front = 0, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b1,     8'b00001010}, // D.10.0, disp_front = 0, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b0,     8'b00000100}, // D.04.0, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b1,     8'b00001100}, // D.12.0, disp_front = 0, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b0,     8'b00000010}, // D.02.0, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b0,     8'b00000001}, // D.01.0, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b0,     8'b00000000}, // D.00.0, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b0,     8'b00000000}, // D.00.0, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b1,     8'b00010001}, // D.17.0, disp_front = 0, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b1,     8'b00010010}, // D.18.0, disp_front = 0, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b0,     8'b00011000}, // D.24.0, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b1,     8'b00010100}, // D.20.0, disp_front = 0, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b0,     8'b00011111}, // D.31.0, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b0,     8'b00010000}, // D.16.0, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b0,     8'b00000000}, // D.00.0, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b1,     8'b00000111}, // D.07.0, disp_front = 0, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b0,     8'b00000000}, // D.00.0, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b0,     8'b00001111}, // D.15.0, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b0,     8'b00000000}, // D.00.0, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b0,     8'b00011100}, // D.28.0, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b0,     8'b00000000}, // D.00.0, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b0,     8'b00000000}, // D.00.0, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b0,     8'b00000000}, // D.00.0, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b0,     8'b11100000}, // D.00.7, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b0,     8'b11100000}, // D.00.7, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b0,     8'b11100000}, // D.00.7, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b0,     8'b11111100}, // D.28.7, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b0,     8'b11100000}, // D.00.7, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b0,     8'b11101111}, // D.15.7, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b0,     8'b11100000}, // D.00.7, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b1,     8'b11100111}, // D.07.7, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b0,     8'b11100000}, // D.00.7, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b0,     8'b11110000}, // D.16.7, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b0,     8'b11111111}, // D.31.7, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b1,     8'b11101011}, // D.11.7, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b0,     8'b11111000}, // D.24.7, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b1,     8'b11101101}, // D.13.7, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b1,     8'b11101110}, // D.14.7, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b0,     1'b1,     1'b0,     1'b0,     8'b11100000}, // D.00.7, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 0
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b0,     8'b11100000}, // D.00.7, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b0,     8'b11100001}, // D.01.7, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b0,     8'b11100010}, // D.02.7, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b1,     8'b11110011}, // D.19.7, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b0,     8'b11100100}, // D.04.7, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b1,     8'b11110101}, // D.21.7, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b1,     8'b11110110}, // D.22.7, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b0,     1'b0,     1'b1,     1'b0,     8'b11110111}, // K.23.7, disp_front = 0, disp_end = 0, K = 1, code_err = 0, disp_err = 0
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b0,     8'b11101000}, // D.08.7, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b1,     8'b11111001}, // D.25.7, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b1,     8'b11111010}, // D.26.7, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b0,     1'b0,     1'b1,     1'b0,     8'b11111011}, // K.27.7, disp_front = 0, disp_end = 0, K = 1, code_err = 0, disp_err = 0
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b1,     8'b11111100}, // D.28.7, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b0,     1'b0,     1'b1,     1'b0,     8'b11111101}, // K.29.7, disp_front = 0, disp_end = 0, K = 1, code_err = 0, disp_err = 0
     {1'b0,       1'b0,     1'b0,     1'b1,     1'b0,     8'b11111110}, // K.30.7, disp_front = 0, disp_end = 0, K = 1, code_err = 0, disp_err = 0
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b0,     8'b11100000}, // D.00.7, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b0,     8'b11100000}, // D.00.7, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b0,     8'b11111110}, // D.30.7, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b0,     8'b11111101}, // D.29.7, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b1,     8'b11100011}, // D.03.7, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b0,     8'b11111011}, // D.27.7, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b1,     8'b11100101}, // D.05.7, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b1,     8'b11100110}, // D.06.7, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b0,     8'b11101000}, // D.08.7, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b0,     8'b11110111}, // D.23.7, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b1,     8'b11101001}, // D.09.7, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b1,     8'b11101010}, // D.10.7, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b0,     8'b11100100}, // D.04.7, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b1,     8'b11101100}, // D.12.7, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b0,     8'b11100010}, // D.02.7, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b0,     8'b11100001}, // D.01.7, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b0,     8'b11100000}, // D.00.7, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b0,     8'b11100000}, // D.00.7, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b1,     8'b11110001}, // D.17.7, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b1,     8'b11110010}, // D.18.7, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b0,     8'b11111000}, // D.24.7, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b1,     8'b11110100}, // D.20.7, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b0,     8'b11111111}, // D.31.7, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b0,     8'b11110000}, // D.16.7, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b0,     8'b11100000}, // D.00.7, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b1,     8'b11100111}, // D.07.7, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b0,     8'b11100000}, // D.00.7, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b0,     8'b11101111}, // D.15.7, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b0,     8'b11100000}, // D.00.7, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b0,     1'b0,     1'b1,     1'b0,     8'b11111100}, // K.28.7, disp_front = 0, disp_end = 0, K = 1, code_err = 0, disp_err = 0
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b0,     8'b11100000}, // D.00.7, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b0,     8'b11100000}, // D.00.7, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b0,     8'b11100000}, // D.00.7, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b0,     8'b00000000}, // D.00.0, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b0,     8'b00000000}, // D.00.0, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b0,     8'b00000000}, // D.00.0, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b0,     8'b00011100}, // D.28.0, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b0,     8'b00000000}, // D.00.0, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b0,     8'b00001111}, // D.15.0, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b0,     8'b00000000}, // D.00.0, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b1,     8'b00000111}, // D.07.0, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b0,     8'b00000000}, // D.00.0, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b0,     8'b00010000}, // D.16.0, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b0,     8'b00011111}, // D.31.0, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b1,     8'b00001011}, // D.11.0, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b0,     8'b00011000}, // D.24.0, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b1,     8'b00001101}, // D.13.0, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b1,     8'b00001110}, // D.14.0, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b0,     1'b1,     1'b0,     1'b0,     8'b00000000}, // D.00.0, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 0
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b0,     8'b00000000}, // D.00.0, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b0,     8'b00000001}, // D.01.0, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b0,     8'b00000010}, // D.02.0, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b1,     8'b00010011}, // D.19.0, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b0,     8'b00000100}, // D.04.0, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b1,     8'b00010101}, // D.21.0, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b1,     8'b00010110}, // D.22.0, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b0,     8'b00010111}, // D.23.0, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b0,     8'b00001000}, // D.08.0, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b1,     8'b00011001}, // D.25.0, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b1,     8'b00011010}, // D.26.0, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b0,     8'b00011011}, // D.27.0, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b1,     8'b00011100}, // D.28.0, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b0,     8'b00011101}, // D.29.0, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b0,     8'b00011110}, // D.30.0, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b0,     8'b00000000}, // D.00.0, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b0,     8'b00000000}, // D.00.0, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b0,     8'b00011110}, // D.30.0, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b0,     8'b00011101}, // D.29.0, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b1,     8'b00000011}, // D.03.0, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b0,     8'b00011011}, // D.27.0, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b1,     8'b00000101}, // D.05.0, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b1,     8'b00000110}, // D.06.0, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b0,     8'b00001000}, // D.08.0, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b0,     8'b00010111}, // D.23.0, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b1,     8'b00001001}, // D.09.0, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b1,     8'b00001010}, // D.10.0, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b0,     8'b00000100}, // D.04.0, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b1,     8'b00001100}, // D.12.0, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b0,     8'b00000010}, // D.02.0, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b0,     8'b00000001}, // D.01.0, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b0,     8'b00000000}, // D.00.0, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b0,     8'b00000000}, // D.00.0, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b1,     8'b00010001}, // D.17.0, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b1,     8'b00010010}, // D.18.0, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b0,     8'b00011000}, // D.24.0, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b1,     8'b00010100}, // D.20.0, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b0,     8'b00011111}, // D.31.0, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b0,     8'b00010000}, // D.16.0, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b0,     8'b00000000}, // D.00.0, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b1,     8'b00000111}, // D.07.0, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b0,     8'b00000000}, // D.00.0, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b0,     8'b00001111}, // D.15.0, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b0,     8'b00000000}, // D.00.0, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b0,     1'b0,     1'b1,     1'b0,     8'b00011100}, // K.28.0, disp_front = 0, disp_end = 0, K = 1, code_err = 0, disp_err = 0
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b0,     8'b00000000}, // D.00.0, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b0,     8'b00000000}, // D.00.0, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b0,     8'b00000000}, // D.00.0, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b1,     8'b01100000}, // D.00.3, disp_front = 0, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b1,     8'b01100000}, // D.00.3, disp_front = 0, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b1,     8'b01100000}, // D.00.3, disp_front = 0, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b1,     1'b1,     8'b01111100}, // K.28.3, disp_front = 0, disp_end = 1, K = 1, code_err = 0, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b1,     8'b01100000}, // D.00.3, disp_front = 0, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b1,     8'b01101111}, // D.15.3, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b1,     8'b01100000}, // D.00.3, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b0,     8'b01100111}, // D.07.3, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b1,     8'b01100000}, // D.00.3, disp_front = 0, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b1,     8'b01110000}, // D.16.3, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b1,     8'b01111111}, // D.31.3, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b0,     8'b01101011}, // D.11.3, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b1,     8'b01111000}, // D.24.3, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b0,     8'b01101101}, // D.13.3, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b0,     8'b01101110}, // D.14.3, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b0,     1'b1,     1'b0,     1'b1,     8'b01100000}, // D.00.3, disp_front = 0, disp_end = 1, K = 0, code_err = 1, disp_err = 0
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b1,     8'b01100000}, // D.00.3, disp_front = 0, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b1,     8'b01100001}, // D.01.3, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b1,     8'b01100010}, // D.02.3, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b0,     8'b01110011}, // D.19.3, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b1,     8'b01100100}, // D.04.3, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b0,     8'b01110101}, // D.21.3, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b0,     8'b01110110}, // D.22.3, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b1,     8'b01110111}, // D.23.3, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b1,     8'b01101000}, // D.08.3, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b0,     8'b01111001}, // D.25.3, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b0,     8'b01111010}, // D.26.3, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b1,     8'b01111011}, // D.27.3, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b0,     8'b01111100}, // D.28.3, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b1,     8'b01111101}, // D.29.3, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b1,     8'b01111110}, // D.30.3, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b1,     8'b01100000}, // D.00.3, disp_front = 0, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b1,     8'b01100000}, // D.00.3, disp_front = 0, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b1,     8'b01111110}, // D.30.3, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b1,     8'b01111101}, // D.29.3, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b0,     8'b01100011}, // D.03.3, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b1,     8'b01111011}, // D.27.3, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b0,     8'b01100101}, // D.05.3, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b0,     8'b01100110}, // D.06.3, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b1,     8'b01101000}, // D.08.3, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b1,     8'b01110111}, // D.23.3, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b0,     8'b01101001}, // D.09.3, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b0,     8'b01101010}, // D.10.3, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b1,     8'b01100100}, // D.04.3, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b0,     8'b01101100}, // D.12.3, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b1,     8'b01100010}, // D.02.3, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b1,     8'b01100001}, // D.01.3, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b1,     8'b01100000}, // D.00.3, disp_front = 0, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b1,     8'b01100000}, // D.00.3, disp_front = 0, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b0,     8'b01110001}, // D.17.3, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b0,     8'b01110010}, // D.18.3, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b1,     8'b01111000}, // D.24.3, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b0,     8'b01110100}, // D.20.3, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b1,     8'b01111111}, // D.31.3, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b1,     8'b01110000}, // D.16.3, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b1,     8'b01100000}, // D.00.3, disp_front = 0, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b0,     8'b01100111}, // D.07.3, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b1,     8'b01100000}, // D.00.3, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b1,     8'b01101111}, // D.15.3, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b1,     8'b01100000}, // D.00.3, disp_front = 0, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b1,     8'b01111100}, // D.28.3, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b1,     8'b01100000}, // D.00.3, disp_front = 0, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b1,     8'b01100000}, // D.00.3, disp_front = 0, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b1,     8'b01100000}, // D.00.3, disp_front = 0, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b0,     8'b10000000}, // D.00.4, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b0,     8'b10000000}, // D.00.4, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b0,     8'b10000000}, // D.00.4, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b0,     8'b10011100}, // D.28.4, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b0,     8'b10000000}, // D.00.4, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b0,     8'b10001111}, // D.15.4, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b0,     8'b10000000}, // D.00.4, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b1,     8'b10000111}, // D.07.4, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b0,     8'b10000000}, // D.00.4, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b0,     8'b10010000}, // D.16.4, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b0,     8'b10011111}, // D.31.4, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b1,     8'b10001011}, // D.11.4, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b0,     8'b10011000}, // D.24.4, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b1,     8'b10001101}, // D.13.4, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b1,     8'b10001110}, // D.14.4, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b0,     1'b1,     1'b0,     1'b0,     8'b10000000}, // D.00.4, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 0
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b0,     8'b10000000}, // D.00.4, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b0,     8'b10000001}, // D.01.4, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b0,     8'b10000010}, // D.02.4, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b1,     8'b10010011}, // D.19.4, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b0,     8'b10000100}, // D.04.4, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b1,     8'b10010101}, // D.21.4, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b1,     8'b10010110}, // D.22.4, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b0,     8'b10010111}, // D.23.4, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b0,     8'b10001000}, // D.08.4, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b1,     8'b10011001}, // D.25.4, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b1,     8'b10011010}, // D.26.4, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b0,     8'b10011011}, // D.27.4, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b1,     8'b10011100}, // D.28.4, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b0,     8'b10011101}, // D.29.4, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b0,     8'b10011110}, // D.30.4, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b0,     8'b10000000}, // D.00.4, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b0,     8'b10000000}, // D.00.4, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b0,     8'b10011110}, // D.30.4, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b0,     8'b10011101}, // D.29.4, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b1,     8'b10000011}, // D.03.4, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b0,     8'b10011011}, // D.27.4, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b1,     8'b10000101}, // D.05.4, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b1,     8'b10000110}, // D.06.4, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b0,     8'b10001000}, // D.08.4, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b0,     8'b10010111}, // D.23.4, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b1,     8'b10001001}, // D.09.4, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b1,     8'b10001010}, // D.10.4, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b0,     8'b10000100}, // D.04.4, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b1,     8'b10001100}, // D.12.4, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b0,     8'b10000010}, // D.02.4, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b0,     8'b10000001}, // D.01.4, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b0,     8'b10000000}, // D.00.4, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b0,     8'b10000000}, // D.00.4, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b1,     8'b10010001}, // D.17.4, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b1,     8'b10010010}, // D.18.4, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b0,     8'b10011000}, // D.24.4, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b1,     8'b10010100}, // D.20.4, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b0,     8'b10011111}, // D.31.4, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b0,     8'b10010000}, // D.16.4, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b0,     8'b10000000}, // D.00.4, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b1,     8'b10000111}, // D.07.4, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b0,     8'b10000000}, // D.00.4, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b0,     8'b10001111}, // D.15.4, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b0,     8'b10000000}, // D.00.4, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b0,     1'b0,     1'b1,     1'b0,     8'b10011100}, // K.28.4, disp_front = 0, disp_end = 0, K = 1, code_err = 0, disp_err = 0
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b0,     8'b10000000}, // D.00.4, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b0,     8'b10000000}, // D.00.4, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b0,     8'b10000000}, // D.00.4, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b1,     8'b10100000}, // D.00.5, disp_front = 0, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b1,     8'b10100000}, // D.00.5, disp_front = 0, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b1,     8'b10100000}, // D.00.5, disp_front = 0, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b1,     1'b1,     8'b10111100}, // K.28.5, disp_front = 0, disp_end = 1, K = 1, code_err = 0, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b1,     8'b10100000}, // D.00.5, disp_front = 0, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b1,     8'b10101111}, // D.15.5, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b1,     8'b10100000}, // D.00.5, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b0,     8'b10100111}, // D.07.5, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b1,     8'b10100000}, // D.00.5, disp_front = 0, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b1,     8'b10110000}, // D.16.5, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b1,     8'b10111111}, // D.31.5, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b0,     8'b10101011}, // D.11.5, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b1,     8'b10111000}, // D.24.5, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b0,     8'b10101101}, // D.13.5, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b0,     8'b10101110}, // D.14.5, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b0,     1'b1,     1'b0,     1'b1,     8'b10100000}, // D.00.5, disp_front = 0, disp_end = 1, K = 0, code_err = 1, disp_err = 0
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b1,     8'b10100000}, // D.00.5, disp_front = 0, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b1,     8'b10100001}, // D.01.5, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b1,     8'b10100010}, // D.02.5, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b0,     8'b10110011}, // D.19.5, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b1,     8'b10100100}, // D.04.5, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b0,     8'b10110101}, // D.21.5, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b0,     8'b10110110}, // D.22.5, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b1,     8'b10110111}, // D.23.5, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b1,     8'b10101000}, // D.08.5, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b0,     8'b10111001}, // D.25.5, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b0,     8'b10111010}, // D.26.5, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b1,     8'b10111011}, // D.27.5, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b0,     8'b10111100}, // D.28.5, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b1,     8'b10111101}, // D.29.5, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b1,     8'b10111110}, // D.30.5, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b1,     8'b10100000}, // D.00.5, disp_front = 0, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b1,     8'b10100000}, // D.00.5, disp_front = 0, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b1,     8'b10111110}, // D.30.5, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b1,     8'b10111101}, // D.29.5, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b0,     8'b10100011}, // D.03.5, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b1,     8'b10111011}, // D.27.5, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b0,     8'b10100101}, // D.05.5, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b0,     8'b10100110}, // D.06.5, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b1,     8'b10101000}, // D.08.5, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b1,     8'b10110111}, // D.23.5, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b0,     8'b10101001}, // D.09.5, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b0,     8'b10101010}, // D.10.5, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b1,     8'b10100100}, // D.04.5, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b0,     8'b10101100}, // D.12.5, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b1,     8'b10100010}, // D.02.5, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b1,     8'b10100001}, // D.01.5, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b1,     8'b10100000}, // D.00.5, disp_front = 0, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b1,     8'b10100000}, // D.00.5, disp_front = 0, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b0,     8'b10110001}, // D.17.5, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b0,     8'b10110010}, // D.18.5, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b1,     8'b10111000}, // D.24.5, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b0,     8'b10110100}, // D.20.5, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b1,     8'b10111111}, // D.31.5, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b1,     8'b10110000}, // D.16.5, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b1,     8'b10100000}, // D.00.5, disp_front = 0, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b0,     8'b10100111}, // D.07.5, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b1,     8'b10100000}, // D.00.5, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b1,     8'b10101111}, // D.15.5, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b1,     8'b10100000}, // D.00.5, disp_front = 0, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b0,     1'b0,     1'b1,     1'b1,     8'b10111100}, // K.28.5, disp_front = 0, disp_end = 1, K = 1, code_err = 0, disp_err = 0
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b1,     8'b10100000}, // D.00.5, disp_front = 0, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b1,     8'b10100000}, // D.00.5, disp_front = 0, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b1,     8'b10100000}, // D.00.5, disp_front = 0, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b1,     8'b11000000}, // D.00.6, disp_front = 0, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b1,     8'b11000000}, // D.00.6, disp_front = 0, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b1,     8'b11000000}, // D.00.6, disp_front = 0, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b1,     1'b1,     8'b11011100}, // K.28.6, disp_front = 0, disp_end = 1, K = 1, code_err = 0, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b1,     8'b11000000}, // D.00.6, disp_front = 0, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b1,     8'b11001111}, // D.15.6, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b1,     8'b11000000}, // D.00.6, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b0,     8'b11000111}, // D.07.6, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b1,     8'b11000000}, // D.00.6, disp_front = 0, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b1,     8'b11010000}, // D.16.6, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b1,     8'b11011111}, // D.31.6, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b0,     8'b11001011}, // D.11.6, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b1,     8'b11011000}, // D.24.6, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b0,     8'b11001101}, // D.13.6, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b0,     8'b11001110}, // D.14.6, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b0,     1'b1,     1'b0,     1'b1,     8'b11000000}, // D.00.6, disp_front = 0, disp_end = 1, K = 0, code_err = 1, disp_err = 0
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b1,     8'b11000000}, // D.00.6, disp_front = 0, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b1,     8'b11000001}, // D.01.6, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b1,     8'b11000010}, // D.02.6, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b0,     8'b11010011}, // D.19.6, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b1,     8'b11000100}, // D.04.6, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b0,     8'b11010101}, // D.21.6, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b0,     8'b11010110}, // D.22.6, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b1,     8'b11010111}, // D.23.6, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b1,     8'b11001000}, // D.08.6, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b0,     8'b11011001}, // D.25.6, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b0,     8'b11011010}, // D.26.6, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b1,     8'b11011011}, // D.27.6, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b0,     8'b11011100}, // D.28.6, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b1,     8'b11011101}, // D.29.6, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b1,     8'b11011110}, // D.30.6, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b1,     8'b11000000}, // D.00.6, disp_front = 0, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b1,     8'b11000000}, // D.00.6, disp_front = 0, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b1,     8'b11011110}, // D.30.6, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b1,     8'b11011101}, // D.29.6, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b0,     8'b11000011}, // D.03.6, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b1,     8'b11011011}, // D.27.6, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b0,     8'b11000101}, // D.05.6, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b0,     8'b11000110}, // D.06.6, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b1,     8'b11001000}, // D.08.6, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b1,     8'b11010111}, // D.23.6, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b0,     8'b11001001}, // D.09.6, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b0,     8'b11001010}, // D.10.6, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b1,     8'b11000100}, // D.04.6, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b0,     8'b11001100}, // D.12.6, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b1,     8'b11000010}, // D.02.6, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b1,     8'b11000001}, // D.01.6, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b1,     8'b11000000}, // D.00.6, disp_front = 0, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b1,     8'b11000000}, // D.00.6, disp_front = 0, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b0,     8'b11010001}, // D.17.6, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b0,     8'b11010010}, // D.18.6, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b1,     8'b11011000}, // D.24.6, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b0,     8'b11010100}, // D.20.6, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b1,     8'b11011111}, // D.31.6, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b1,     8'b11010000}, // D.16.6, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b1,     8'b11000000}, // D.00.6, disp_front = 0, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b0,     8'b11000111}, // D.07.6, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b1,     8'b11000000}, // D.00.6, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b1,     8'b11001111}, // D.15.6, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b1,     8'b11000000}, // D.00.6, disp_front = 0, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b0,     1'b0,     1'b1,     1'b1,     8'b11011100}, // K.28.6, disp_front = 0, disp_end = 1, K = 1, code_err = 0, disp_err = 0
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b1,     8'b11000000}, // D.00.6, disp_front = 0, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b1,     8'b11000000}, // D.00.6, disp_front = 0, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b1,     8'b11000000}, // D.00.6, disp_front = 0, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b0,     8'b11100000}, // D.00.7, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b0,     8'b11100000}, // D.00.7, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b0,     8'b11100000}, // D.00.7, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b0,     8'b11111100}, // D.28.7, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b0,     8'b11100000}, // D.00.7, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b0,     8'b11101111}, // D.15.7, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b0,     8'b11100000}, // D.00.7, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b1,     8'b11100111}, // D.07.7, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b0,     8'b11100000}, // D.00.7, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b0,     8'b11110000}, // D.16.7, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b0,     8'b11111111}, // D.31.7, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b1,     8'b11101011}, // D.11.7, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b0,     8'b11111000}, // D.24.7, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b1,     8'b11101101}, // D.13.7, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b1,     8'b11101110}, // D.14.7, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b0,     8'b11100000}, // D.00.7, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b0,     8'b11100000}, // D.00.7, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b0,     8'b11100001}, // D.01.7, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b0,     8'b11100010}, // D.02.7, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b1,     8'b11110011}, // D.19.7, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b0,     8'b11100100}, // D.04.7, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b1,     8'b11110101}, // D.21.7, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b1,     8'b11110110}, // D.22.7, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b0,     8'b11110111}, // D.23.7, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b0,     8'b11101000}, // D.08.7, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b1,     8'b11111001}, // D.25.7, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b1,     8'b11111010}, // D.26.7, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b0,     8'b11111011}, // D.27.7, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b1,     8'b11111100}, // D.28.7, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b0,     8'b11111101}, // D.29.7, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b0,     8'b11111110}, // D.30.7, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b0,     8'b11100000}, // D.00.7, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b0,     8'b11100000}, // D.00.7, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b0,     8'b11111110}, // D.30.7, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b0,     8'b11111101}, // D.29.7, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b1,     8'b11100011}, // D.03.7, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b0,     8'b11111011}, // D.27.7, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b1,     8'b11100101}, // D.05.7, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b1,     8'b11100110}, // D.06.7, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b0,     8'b11101000}, // D.08.7, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b0,     8'b11110111}, // D.23.7, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b1,     8'b11101001}, // D.09.7, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b1,     8'b11101010}, // D.10.7, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b0,     8'b11100100}, // D.04.7, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b1,     8'b11101100}, // D.12.7, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b0,     8'b11100010}, // D.02.7, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b0,     8'b11100001}, // D.01.7, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b0,     8'b11100000}, // D.00.7, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b0,     8'b11100000}, // D.00.7, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b1,     8'b11110001}, // D.17.7, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b1,     8'b11110010}, // D.18.7, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b0,     8'b11111000}, // D.24.7, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b1,     8'b11110100}, // D.20.7, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b0,     8'b11111111}, // D.31.7, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b0,     8'b11110000}, // D.16.7, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b0,     8'b11100000}, // D.00.7, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b1,     8'b11100111}, // D.07.7, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b0,     8'b11100000}, // D.00.7, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b0,     8'b11101111}, // D.15.7, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b0,     8'b11100000}, // D.00.7, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b0,     8'b11111100}, // D.28.7, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b0,     8'b11100000}, // D.00.7, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b0,     8'b11100000}, // D.00.7, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b0,     8'b11100000}, // D.00.7, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b0,     8'b11100000}, // D.00.7, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b0,     8'b11100000}, // D.00.7, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b0,     8'b11100000}, // D.00.7, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b0,     8'b11111100}, // D.28.7, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b0,     8'b11100000}, // D.00.7, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b0,     8'b11101111}, // D.15.7, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b0,     8'b11100000}, // D.00.7, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b1,     8'b11100111}, // D.07.7, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b0,     8'b11100000}, // D.00.7, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b0,     8'b11110000}, // D.16.7, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b0,     8'b11111111}, // D.31.7, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b1,     8'b11101011}, // D.11.7, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b0,     8'b11111000}, // D.24.7, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b1,     8'b11101101}, // D.13.7, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b1,     8'b11101110}, // D.14.7, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b0,     1'b1,     1'b0,     1'b0,     8'b11100000}, // D.00.7, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 0
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b0,     8'b11100000}, // D.00.7, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b0,     8'b11100001}, // D.01.7, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b0,     8'b11100010}, // D.02.7, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b1,     8'b11110011}, // D.19.7, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b0,     8'b11100100}, // D.04.7, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b1,     8'b11110101}, // D.21.7, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b1,     8'b11110110}, // D.22.7, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b0,     8'b11110111}, // D.23.7, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b0,     8'b11101000}, // D.08.7, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b1,     8'b11111001}, // D.25.7, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b1,     8'b11111010}, // D.26.7, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b0,     8'b11111011}, // D.27.7, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b1,     8'b11111100}, // D.28.7, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b0,     8'b11111101}, // D.29.7, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b0,     8'b11111110}, // D.30.7, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b0,     8'b11100000}, // D.00.7, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b0,     8'b11100000}, // D.00.7, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b0,     8'b11111110}, // D.30.7, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b0,     8'b11111101}, // D.29.7, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b1,     8'b11100011}, // D.03.7, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b0,     8'b11111011}, // D.27.7, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b1,     8'b11100101}, // D.05.7, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b1,     8'b11100110}, // D.06.7, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b0,     8'b11101000}, // D.08.7, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b0,     8'b11110111}, // D.23.7, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b1,     8'b11101001}, // D.09.7, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b1,     8'b11101010}, // D.10.7, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b0,     8'b11100100}, // D.04.7, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b1,     8'b11101100}, // D.12.7, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b0,     8'b11100010}, // D.02.7, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b0,     8'b11100001}, // D.01.7, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b0,     8'b11100000}, // D.00.7, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b0,     8'b11100000}, // D.00.7, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b1,     8'b11110001}, // D.17.7, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b1,     8'b11110010}, // D.18.7, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b0,     8'b11111000}, // D.24.7, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b1,     8'b11110100}, // D.20.7, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b0,     8'b11111111}, // D.31.7, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b0,     8'b11110000}, // D.16.7, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b0,     8'b11100000}, // D.00.7, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b1,     8'b11100111}, // D.07.7, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b0,     8'b11100000}, // D.00.7, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b0,     8'b11101111}, // D.15.7, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b0,     8'b11100000}, // D.00.7, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b0,     8'b11111100}, // D.28.7, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b0,     8'b11100000}, // D.00.7, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b0,     8'b11100000}, // D.00.7, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b0,     8'b11100000}, // D.00.7, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b1,     8'b00100000}, // D.00.1, disp_front = 0, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b1,     8'b00100000}, // D.00.1, disp_front = 0, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b1,     8'b00100000}, // D.00.1, disp_front = 0, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b1,     1'b1,     8'b00111100}, // K.28.1, disp_front = 0, disp_end = 1, K = 1, code_err = 0, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b1,     8'b00100000}, // D.00.1, disp_front = 0, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b1,     8'b00101111}, // D.15.1, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b1,     8'b00100000}, // D.00.1, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b0,     8'b00100111}, // D.07.1, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b1,     8'b00100000}, // D.00.1, disp_front = 0, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b1,     8'b00110000}, // D.16.1, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b1,     8'b00111111}, // D.31.1, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b0,     8'b00101011}, // D.11.1, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b1,     8'b00111000}, // D.24.1, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b0,     8'b00101101}, // D.13.1, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b0,     8'b00101110}, // D.14.1, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b0,     1'b1,     1'b0,     1'b1,     8'b00100000}, // D.00.1, disp_front = 0, disp_end = 1, K = 0, code_err = 1, disp_err = 0
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b1,     8'b00100000}, // D.00.1, disp_front = 0, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b1,     8'b00100001}, // D.01.1, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b1,     8'b00100010}, // D.02.1, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b0,     8'b00110011}, // D.19.1, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b1,     8'b00100100}, // D.04.1, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b0,     8'b00110101}, // D.21.1, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b0,     8'b00110110}, // D.22.1, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b1,     8'b00110111}, // D.23.1, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b1,     8'b00101000}, // D.08.1, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b0,     8'b00111001}, // D.25.1, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b0,     8'b00111010}, // D.26.1, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b1,     8'b00111011}, // D.27.1, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b0,     8'b00111100}, // D.28.1, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b1,     8'b00111101}, // D.29.1, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b1,     8'b00111110}, // D.30.1, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b1,     8'b00100000}, // D.00.1, disp_front = 0, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b1,     8'b00100000}, // D.00.1, disp_front = 0, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b1,     8'b00111110}, // D.30.1, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b1,     8'b00111101}, // D.29.1, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b0,     8'b00100011}, // D.03.1, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b1,     8'b00111011}, // D.27.1, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b0,     8'b00100101}, // D.05.1, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b0,     8'b00100110}, // D.06.1, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b1,     8'b00101000}, // D.08.1, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b1,     8'b00110111}, // D.23.1, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b0,     8'b00101001}, // D.09.1, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b0,     8'b00101010}, // D.10.1, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b1,     8'b00100100}, // D.04.1, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b0,     8'b00101100}, // D.12.1, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b1,     8'b00100010}, // D.02.1, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b1,     8'b00100001}, // D.01.1, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b1,     8'b00100000}, // D.00.1, disp_front = 0, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b1,     8'b00100000}, // D.00.1, disp_front = 0, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b0,     8'b00110001}, // D.17.1, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b0,     8'b00110010}, // D.18.1, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b1,     8'b00111000}, // D.24.1, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b0,     8'b00110100}, // D.20.1, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b1,     8'b00111111}, // D.31.1, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b1,     8'b00110000}, // D.16.1, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b1,     8'b00100000}, // D.00.1, disp_front = 0, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b0,     8'b00100111}, // D.07.1, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b1,     8'b00100000}, // D.00.1, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b1,     8'b00101111}, // D.15.1, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b1,     8'b00100000}, // D.00.1, disp_front = 0, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b0,     1'b0,     1'b1,     1'b1,     8'b00111100}, // K.28.1, disp_front = 0, disp_end = 1, K = 1, code_err = 0, disp_err = 0
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b1,     8'b00100000}, // D.00.1, disp_front = 0, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b1,     8'b00100000}, // D.00.1, disp_front = 0, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b1,     8'b00100000}, // D.00.1, disp_front = 0, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b1,     8'b01000000}, // D.00.2, disp_front = 0, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b1,     8'b01000000}, // D.00.2, disp_front = 0, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b1,     8'b01000000}, // D.00.2, disp_front = 0, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b1,     1'b1,     8'b01011100}, // K.28.2, disp_front = 0, disp_end = 1, K = 1, code_err = 0, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b1,     8'b01000000}, // D.00.2, disp_front = 0, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b1,     8'b01001111}, // D.15.2, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b1,     8'b01000000}, // D.00.2, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b0,     8'b01000111}, // D.07.2, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b1,     8'b01000000}, // D.00.2, disp_front = 0, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b1,     8'b01010000}, // D.16.2, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b1,     8'b01011111}, // D.31.2, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b0,     8'b01001011}, // D.11.2, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b1,     8'b01011000}, // D.24.2, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b0,     8'b01001101}, // D.13.2, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b0,     8'b01001110}, // D.14.2, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b0,     1'b1,     1'b0,     1'b1,     8'b01000000}, // D.00.2, disp_front = 0, disp_end = 1, K = 0, code_err = 1, disp_err = 0
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b1,     8'b01000000}, // D.00.2, disp_front = 0, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b1,     8'b01000001}, // D.01.2, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b1,     8'b01000010}, // D.02.2, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b0,     8'b01010011}, // D.19.2, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b1,     8'b01000100}, // D.04.2, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b0,     8'b01010101}, // D.21.2, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b0,     8'b01010110}, // D.22.2, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b1,     8'b01010111}, // D.23.2, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b1,     8'b01001000}, // D.08.2, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b0,     8'b01011001}, // D.25.2, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b0,     8'b01011010}, // D.26.2, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b1,     8'b01011011}, // D.27.2, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b0,     8'b01011100}, // D.28.2, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b1,     8'b01011101}, // D.29.2, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b1,     8'b01011110}, // D.30.2, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b1,     8'b01000000}, // D.00.2, disp_front = 0, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b1,     8'b01000000}, // D.00.2, disp_front = 0, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b1,     8'b01011110}, // D.30.2, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b1,     8'b01011101}, // D.29.2, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b0,     8'b01000011}, // D.03.2, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b1,     8'b01011011}, // D.27.2, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b0,     8'b01000101}, // D.05.2, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b0,     8'b01000110}, // D.06.2, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b1,     8'b01001000}, // D.08.2, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b1,     8'b01010111}, // D.23.2, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b0,     8'b01001001}, // D.09.2, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b0,     8'b01001010}, // D.10.2, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b1,     8'b01000100}, // D.04.2, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b0,     8'b01001100}, // D.12.2, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b1,     8'b01000010}, // D.02.2, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b1,     8'b01000001}, // D.01.2, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b1,     8'b01000000}, // D.00.2, disp_front = 0, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b1,     8'b01000000}, // D.00.2, disp_front = 0, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b0,     8'b01010001}, // D.17.2, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b0,     8'b01010010}, // D.18.2, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b1,     8'b01011000}, // D.24.2, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b0,     8'b01010100}, // D.20.2, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b1,     8'b01011111}, // D.31.2, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b1,     8'b01010000}, // D.16.2, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b1,     8'b01000000}, // D.00.2, disp_front = 0, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b0,     8'b01000111}, // D.07.2, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b1,     8'b01000000}, // D.00.2, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b1,     8'b01001111}, // D.15.2, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b1,     8'b01000000}, // D.00.2, disp_front = 0, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b0,     1'b0,     1'b1,     1'b1,     8'b01011100}, // K.28.2, disp_front = 0, disp_end = 1, K = 1, code_err = 0, disp_err = 0
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b1,     8'b01000000}, // D.00.2, disp_front = 0, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b1,     8'b01000000}, // D.00.2, disp_front = 0, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b1,     8'b01000000}, // D.00.2, disp_front = 0, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b0,     8'b10000000}, // D.00.4, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b0,     8'b10000000}, // D.00.4, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b0,     8'b10000000}, // D.00.4, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b1,     1'b0,     8'b10011100}, // K.28.4, disp_front = 0, disp_end = 0, K = 1, code_err = 0, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b0,     8'b10000000}, // D.00.4, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b0,     8'b10001111}, // D.15.4, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b0,     8'b10000000}, // D.00.4, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b1,     8'b10000111}, // D.07.4, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b0,     8'b10000000}, // D.00.4, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b0,     8'b10010000}, // D.16.4, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b0,     8'b10011111}, // D.31.4, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b1,     8'b10001011}, // D.11.4, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b0,     8'b10011000}, // D.24.4, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b1,     8'b10001101}, // D.13.4, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b1,     8'b10001110}, // D.14.4, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b0,     8'b10000000}, // D.00.4, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b0,     8'b10000000}, // D.00.4, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b0,     8'b10000001}, // D.01.4, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b0,     8'b10000010}, // D.02.4, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b1,     8'b10010011}, // D.19.4, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b0,     8'b10000100}, // D.04.4, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b1,     8'b10010101}, // D.21.4, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b1,     8'b10010110}, // D.22.4, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b0,     8'b10010111}, // D.23.4, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b0,     8'b10001000}, // D.08.4, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b1,     8'b10011001}, // D.25.4, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b1,     8'b10011010}, // D.26.4, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b0,     8'b10011011}, // D.27.4, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b1,     8'b10011100}, // D.28.4, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b0,     8'b10011101}, // D.29.4, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b0,     8'b10011110}, // D.30.4, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b0,     8'b10000000}, // D.00.4, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b0,     8'b10000000}, // D.00.4, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b0,     8'b10011110}, // D.30.4, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b0,     8'b10011101}, // D.29.4, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b1,     8'b10000011}, // D.03.4, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b0,     8'b10011011}, // D.27.4, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b1,     8'b10000101}, // D.05.4, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b1,     8'b10000110}, // D.06.4, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b0,     8'b10001000}, // D.08.4, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b0,     8'b10010111}, // D.23.4, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b1,     8'b10001001}, // D.09.4, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b1,     8'b10001010}, // D.10.4, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b0,     8'b10000100}, // D.04.4, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b1,     8'b10001100}, // D.12.4, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b0,     8'b10000010}, // D.02.4, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b0,     8'b10000001}, // D.01.4, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b0,     8'b10000000}, // D.00.4, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b0,     8'b10000000}, // D.00.4, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b1,     8'b10010001}, // D.17.4, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b1,     8'b10010010}, // D.18.4, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b0,     8'b10011000}, // D.24.4, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b1,     8'b10010100}, // D.20.4, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b0,     8'b10011111}, // D.31.4, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b0,     8'b10010000}, // D.16.4, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b0,     8'b10000000}, // D.00.4, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b1,     8'b10000111}, // D.07.4, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b0,     8'b10000000}, // D.00.4, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b0,     8'b10001111}, // D.15.4, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b0,     8'b10000000}, // D.00.4, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b0,     8'b10011100}, // D.28.4, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b0,     8'b10000000}, // D.00.4, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b0,     8'b10000000}, // D.00.4, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b0,     8'b10000000}, // D.00.4, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b1,     8'b01100000}, // D.00.3, disp_front = 0, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b1,     8'b01100000}, // D.00.3, disp_front = 0, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b1,     8'b01100000}, // D.00.3, disp_front = 0, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b1,     8'b01111100}, // D.28.3, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b1,     8'b01100000}, // D.00.3, disp_front = 0, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b1,     8'b01101111}, // D.15.3, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b1,     8'b01100000}, // D.00.3, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b0,     8'b01100111}, // D.07.3, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b1,     8'b01100000}, // D.00.3, disp_front = 0, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b1,     8'b01110000}, // D.16.3, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b1,     8'b01111111}, // D.31.3, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b0,     8'b01101011}, // D.11.3, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b1,     8'b01111000}, // D.24.3, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b0,     8'b01101101}, // D.13.3, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b0,     8'b01101110}, // D.14.3, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b0,     1'b1,     1'b0,     1'b1,     8'b01100000}, // D.00.3, disp_front = 0, disp_end = 1, K = 0, code_err = 1, disp_err = 0
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b1,     8'b01100000}, // D.00.3, disp_front = 0, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b1,     8'b01100001}, // D.01.3, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b1,     8'b01100010}, // D.02.3, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b0,     8'b01110011}, // D.19.3, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b1,     8'b01100100}, // D.04.3, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b0,     8'b01110101}, // D.21.3, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b0,     8'b01110110}, // D.22.3, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b1,     8'b01110111}, // D.23.3, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b1,     8'b01101000}, // D.08.3, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b0,     8'b01111001}, // D.25.3, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b0,     8'b01111010}, // D.26.3, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b1,     8'b01111011}, // D.27.3, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b0,     8'b01111100}, // D.28.3, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b1,     8'b01111101}, // D.29.3, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b1,     8'b01111110}, // D.30.3, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b1,     8'b01100000}, // D.00.3, disp_front = 0, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b1,     8'b01100000}, // D.00.3, disp_front = 0, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b1,     8'b01111110}, // D.30.3, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b1,     8'b01111101}, // D.29.3, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b0,     8'b01100011}, // D.03.3, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b1,     8'b01111011}, // D.27.3, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b0,     8'b01100101}, // D.05.3, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b0,     8'b01100110}, // D.06.3, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b1,     8'b01101000}, // D.08.3, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b1,     8'b01110111}, // D.23.3, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b0,     8'b01101001}, // D.09.3, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b0,     8'b01101010}, // D.10.3, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b1,     8'b01100100}, // D.04.3, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b0,     8'b01101100}, // D.12.3, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b1,     8'b01100010}, // D.02.3, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b1,     8'b01100001}, // D.01.3, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b1,     8'b01100000}, // D.00.3, disp_front = 0, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b1,     8'b01100000}, // D.00.3, disp_front = 0, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b0,     8'b01110001}, // D.17.3, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b0,     8'b01110010}, // D.18.3, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b1,     8'b01111000}, // D.24.3, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b0,     8'b01110100}, // D.20.3, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b1,     8'b01111111}, // D.31.3, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b1,     8'b01110000}, // D.16.3, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b1,     8'b01100000}, // D.00.3, disp_front = 0, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b0,     8'b01100111}, // D.07.3, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b1,     8'b01100000}, // D.00.3, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b1,     8'b01101111}, // D.15.3, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b1,     8'b01100000}, // D.00.3, disp_front = 0, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b0,     1'b0,     1'b1,     1'b1,     8'b01111100}, // K.28.3, disp_front = 0, disp_end = 1, K = 1, code_err = 0, disp_err = 0
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b1,     8'b01100000}, // D.00.3, disp_front = 0, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b1,     8'b01100000}, // D.00.3, disp_front = 0, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b1,     8'b01100000}, // D.00.3, disp_front = 0, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b0,     8'b00000000}, // D.00.0, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b0,     8'b00000000}, // D.00.0, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b0,     8'b00000000}, // D.00.0, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b1,     1'b0,     8'b00011100}, // K.28.0, disp_front = 0, disp_end = 0, K = 1, code_err = 0, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b0,     8'b00000000}, // D.00.0, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b0,     8'b00001111}, // D.15.0, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b0,     8'b00000000}, // D.00.0, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b1,     8'b00000111}, // D.07.0, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b0,     8'b00000000}, // D.00.0, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b0,     8'b00010000}, // D.16.0, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b0,     8'b00011111}, // D.31.0, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b1,     8'b00001011}, // D.11.0, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b0,     8'b00011000}, // D.24.0, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b1,     8'b00001101}, // D.13.0, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b1,     8'b00001110}, // D.14.0, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b0,     8'b00000000}, // D.00.0, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b0,     8'b00000000}, // D.00.0, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b0,     8'b00000001}, // D.01.0, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b0,     8'b00000010}, // D.02.0, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b1,     8'b00010011}, // D.19.0, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b0,     8'b00000100}, // D.04.0, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b1,     8'b00010101}, // D.21.0, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b1,     8'b00010110}, // D.22.0, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b0,     8'b00010111}, // D.23.0, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b0,     8'b00001000}, // D.08.0, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b1,     8'b00011001}, // D.25.0, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b1,     8'b00011010}, // D.26.0, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b0,     8'b00011011}, // D.27.0, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b1,     8'b00011100}, // D.28.0, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b0,     8'b00011101}, // D.29.0, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b0,     8'b00011110}, // D.30.0, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b0,     8'b00000000}, // D.00.0, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b0,     8'b00000000}, // D.00.0, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b0,     8'b00011110}, // D.30.0, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b0,     8'b00011101}, // D.29.0, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b1,     8'b00000011}, // D.03.0, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b0,     8'b00011011}, // D.27.0, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b1,     8'b00000101}, // D.05.0, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b1,     8'b00000110}, // D.06.0, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b0,     8'b00001000}, // D.08.0, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b0,     8'b00010111}, // D.23.0, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b1,     8'b00001001}, // D.09.0, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b1,     8'b00001010}, // D.10.0, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b0,     8'b00000100}, // D.04.0, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b1,     8'b00001100}, // D.12.0, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b0,     8'b00000010}, // D.02.0, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b0,     8'b00000001}, // D.01.0, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b0,     8'b00000000}, // D.00.0, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b0,     8'b00000000}, // D.00.0, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b1,     8'b00010001}, // D.17.0, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b1,     8'b00010010}, // D.18.0, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b0,     8'b00011000}, // D.24.0, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b1,     8'b00010100}, // D.20.0, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b0,     8'b00011111}, // D.31.0, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b0,     8'b00010000}, // D.16.0, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b0,     8'b00000000}, // D.00.0, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b1,     8'b00000111}, // D.07.0, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b0,     8'b00000000}, // D.00.0, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b0,     8'b00001111}, // D.15.0, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b0,     8'b00000000}, // D.00.0, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b0,     8'b00011100}, // D.28.0, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b0,     8'b00000000}, // D.00.0, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b0,     8'b00000000}, // D.00.0, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b0,     8'b00000000}, // D.00.0, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b0,     8'b11100000}, // D.00.7, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b0,     8'b11100000}, // D.00.7, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b0,     8'b11100000}, // D.00.7, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b1,     1'b0,     8'b11111100}, // K.28.7, disp_front = 0, disp_end = 0, K = 1, code_err = 0, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b0,     8'b11100000}, // D.00.7, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b0,     8'b11101111}, // D.15.7, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b0,     8'b11100000}, // D.00.7, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b1,     8'b11100111}, // D.07.7, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b0,     8'b11100000}, // D.00.7, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b0,     8'b11110000}, // D.16.7, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b0,     8'b11111111}, // D.31.7, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b1,     8'b11101011}, // D.11.7, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b0,     8'b11111000}, // D.24.7, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b1,     8'b11101101}, // D.13.7, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b1,     8'b11101110}, // D.14.7, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b0,     8'b11100000}, // D.00.7, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b0,     8'b11100000}, // D.00.7, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b0,     8'b11100001}, // D.01.7, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b0,     8'b11100010}, // D.02.7, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b1,     8'b11110011}, // D.19.7, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b0,     8'b11100100}, // D.04.7, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b1,     8'b11110101}, // D.21.7, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b1,     8'b11110110}, // D.22.7, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b0,     8'b11110111}, // D.23.7, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b0,     8'b11101000}, // D.08.7, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b1,     8'b11111001}, // D.25.7, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b1,     8'b11111010}, // D.26.7, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b0,     8'b11111011}, // D.27.7, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b1,     8'b11111100}, // D.28.7, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b0,     8'b11111101}, // D.29.7, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b0,     8'b11111110}, // D.30.7, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b0,     8'b11100000}, // D.00.7, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b0,     8'b11100000}, // D.00.7, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b1,     1'b0,     8'b11111110}, // K.30.7, disp_front = 0, disp_end = 0, K = 1, code_err = 0, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b1,     1'b0,     8'b11111101}, // K.29.7, disp_front = 0, disp_end = 0, K = 1, code_err = 0, disp_err = 1
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b1,     8'b11100011}, // D.03.7, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b1,     1'b0,     1'b1,     1'b0,     8'b11111011}, // K.27.7, disp_front = 0, disp_end = 0, K = 1, code_err = 0, disp_err = 1
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b1,     8'b11100101}, // D.05.7, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b1,     8'b11100110}, // D.06.7, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b0,     8'b11101000}, // D.08.7, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b1,     1'b0,     8'b11110111}, // K.23.7, disp_front = 0, disp_end = 0, K = 1, code_err = 0, disp_err = 1
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b1,     8'b11101001}, // D.09.7, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b1,     8'b11101010}, // D.10.7, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b0,     8'b11100100}, // D.04.7, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b1,     8'b11101100}, // D.12.7, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b0,     8'b11100010}, // D.02.7, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b0,     8'b11100001}, // D.01.7, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b0,     8'b11100000}, // D.00.7, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b0,     8'b11100000}, // D.00.7, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b1,     8'b11110001}, // D.17.7, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b1,     8'b11110010}, // D.18.7, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b0,     8'b11111000}, // D.24.7, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b1,     8'b11110100}, // D.20.7, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b0,     8'b11111111}, // D.31.7, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b0,     8'b11110000}, // D.16.7, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b0,     8'b11100000}, // D.00.7, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b0,     1'b0,     1'b0,     1'b1,     8'b11100111}, // D.07.7, disp_front = 0, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b0,     8'b11100000}, // D.00.7, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b0,     8'b11101111}, // D.15.7, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b0,     8'b11100000}, // D.00.7, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b0,     1'b0,     1'b0,     8'b11111100}, // D.28.7, disp_front = 0, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b0,     8'b11100000}, // D.00.7, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b0,     8'b11100000}, // D.00.7, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b0,     8'b11100000}, // D.00.7, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b0,     8'b00000000}, // D.00.0, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b0,     8'b00000000}, // D.00.0, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b0,     8'b00000000}, // D.00.0, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b0,     8'b00011100}, // D.28.0, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b0,     8'b00000000}, // D.00.0, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b0,     8'b00001111}, // D.15.0, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b0,     8'b00000000}, // D.00.0, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b1,     8'b00000111}, // D.07.0, disp_front = 0, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b0,     8'b00000000}, // D.00.0, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b0,     8'b00010000}, // D.16.0, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b0,     8'b00011111}, // D.31.0, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b1,     8'b00001011}, // D.11.0, disp_front = 0, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b0,     8'b00011000}, // D.24.0, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b1,     8'b00001101}, // D.13.0, disp_front = 0, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b1,     8'b00001110}, // D.14.0, disp_front = 0, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b0,     8'b00000000}, // D.00.0, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b0,     8'b00000000}, // D.00.0, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b0,     8'b00000001}, // D.01.0, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b0,     8'b00000010}, // D.02.0, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b1,     8'b00010011}, // D.19.0, disp_front = 0, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b0,     8'b00000100}, // D.04.0, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b1,     8'b00010101}, // D.21.0, disp_front = 0, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b1,     8'b00010110}, // D.22.0, disp_front = 0, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b0,     8'b00010111}, // D.23.0, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b0,     8'b00001000}, // D.08.0, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b1,     8'b00011001}, // D.25.0, disp_front = 0, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b1,     8'b00011010}, // D.26.0, disp_front = 0, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b0,     8'b00011011}, // D.27.0, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b1,     8'b00011100}, // D.28.0, disp_front = 0, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b0,     8'b00011101}, // D.29.0, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b0,     8'b00011110}, // D.30.0, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b0,     8'b00000000}, // D.00.0, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b0,     8'b00000000}, // D.00.0, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b0,     8'b00011110}, // D.30.0, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b0,     8'b00011101}, // D.29.0, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b1,     8'b00000011}, // D.03.0, disp_front = 0, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b0,     8'b00011011}, // D.27.0, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b1,     8'b00000101}, // D.05.0, disp_front = 0, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b1,     8'b00000110}, // D.06.0, disp_front = 0, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b0,     8'b00001000}, // D.08.0, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b0,     8'b00010111}, // D.23.0, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b1,     8'b00001001}, // D.09.0, disp_front = 0, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b1,     8'b00001010}, // D.10.0, disp_front = 0, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b0,     8'b00000100}, // D.04.0, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b1,     8'b00001100}, // D.12.0, disp_front = 0, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b0,     8'b00000010}, // D.02.0, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b0,     8'b00000001}, // D.01.0, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b0,     8'b00000000}, // D.00.0, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b0,     8'b00000000}, // D.00.0, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b1,     8'b00010001}, // D.17.0, disp_front = 0, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b1,     8'b00010010}, // D.18.0, disp_front = 0, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b0,     8'b00011000}, // D.24.0, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b1,     8'b00010100}, // D.20.0, disp_front = 0, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b0,     8'b00011111}, // D.31.0, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b0,     8'b00010000}, // D.16.0, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b0,     8'b00000000}, // D.00.0, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b1,     8'b00000111}, // D.07.0, disp_front = 0, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b0,     8'b00000000}, // D.00.0, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b0,     8'b00001111}, // D.15.0, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b0,     8'b00000000}, // D.00.0, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b0,     8'b00011100}, // D.28.0, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b0,     8'b00000000}, // D.00.0, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b0,     8'b00000000}, // D.00.0, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b0,       1'b1,     1'b1,     1'b0,     1'b0,     8'b00000000}, // D.00.0, disp_front = 0, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b1,     8'b00000000}, // D.00.0, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b1,     8'b00000000}, // D.00.0, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b1,     8'b00000000}, // D.00.0, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b1,     8'b00011100}, // D.28.0, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b1,     8'b00000000}, // D.00.0, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b1,     8'b00001111}, // D.15.0, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b1,     8'b00000000}, // D.00.0, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b0,     8'b00000111}, // D.07.0, disp_front = 1, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b1,     8'b00000000}, // D.00.0, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b1,     8'b00010000}, // D.16.0, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b1,     8'b00011111}, // D.31.0, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b0,     8'b00001011}, // D.11.0, disp_front = 1, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b1,     8'b00011000}, // D.24.0, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b0,     8'b00001101}, // D.13.0, disp_front = 1, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b0,     8'b00001110}, // D.14.0, disp_front = 1, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b1,     8'b00000000}, // D.00.0, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b1,     8'b00000000}, // D.00.0, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b1,     8'b00000001}, // D.01.0, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b1,     8'b00000010}, // D.02.0, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b0,     8'b00010011}, // D.19.0, disp_front = 1, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b1,     8'b00000100}, // D.04.0, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b0,     8'b00010101}, // D.21.0, disp_front = 1, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b0,     8'b00010110}, // D.22.0, disp_front = 1, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b1,     8'b00010111}, // D.23.0, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b1,     8'b00001000}, // D.08.0, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b0,     8'b00011001}, // D.25.0, disp_front = 1, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b0,     8'b00011010}, // D.26.0, disp_front = 1, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b1,     8'b00011011}, // D.27.0, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b0,     8'b00011100}, // D.28.0, disp_front = 1, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b1,     8'b00011101}, // D.29.0, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b1,     8'b00011110}, // D.30.0, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b1,     8'b00000000}, // D.00.0, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b1,     8'b00000000}, // D.00.0, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b1,     8'b00011110}, // D.30.0, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b1,     8'b00011101}, // D.29.0, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b0,     8'b00000011}, // D.03.0, disp_front = 1, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b1,     8'b00011011}, // D.27.0, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b0,     8'b00000101}, // D.05.0, disp_front = 1, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b0,     8'b00000110}, // D.06.0, disp_front = 1, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b1,     8'b00001000}, // D.08.0, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b1,     8'b00010111}, // D.23.0, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b0,     8'b00001001}, // D.09.0, disp_front = 1, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b0,     8'b00001010}, // D.10.0, disp_front = 1, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b1,     8'b00000100}, // D.04.0, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b0,     8'b00001100}, // D.12.0, disp_front = 1, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b1,     8'b00000010}, // D.02.0, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b1,     8'b00000001}, // D.01.0, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b1,     8'b00000000}, // D.00.0, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b1,     8'b00000000}, // D.00.0, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b0,     8'b00010001}, // D.17.0, disp_front = 1, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b0,     8'b00010010}, // D.18.0, disp_front = 1, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b1,     8'b00011000}, // D.24.0, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b0,     8'b00010100}, // D.20.0, disp_front = 1, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b1,     8'b00011111}, // D.31.0, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b1,     8'b00010000}, // D.16.0, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b1,     8'b00000000}, // D.00.0, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b0,     8'b00000111}, // D.07.0, disp_front = 1, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b1,     8'b00000000}, // D.00.0, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b1,     8'b00001111}, // D.15.0, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b1,     8'b00000000}, // D.00.0, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b1,     8'b00011100}, // D.28.0, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b1,     8'b00000000}, // D.00.0, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b1,     8'b00000000}, // D.00.0, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b1,     8'b00000000}, // D.00.0, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b1,     8'b11100000}, // D.00.7, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b1,     8'b11100000}, // D.00.7, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b1,     8'b11100000}, // D.00.7, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b1,     8'b11111100}, // D.28.7, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b1,     8'b11100000}, // D.00.7, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b1,     8'b11101111}, // D.15.7, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b1,     8'b11100000}, // D.00.7, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b0,     8'b11100111}, // D.07.7, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b1,     8'b11100000}, // D.00.7, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b1,     8'b11110000}, // D.16.7, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b1,     8'b11111111}, // D.31.7, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b0,     8'b11101011}, // D.11.7, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b1,     8'b11111000}, // D.24.7, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b0,     8'b11101101}, // D.13.7, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b0,     8'b11101110}, // D.14.7, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b1,     8'b11100000}, // D.00.7, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b1,     8'b11100000}, // D.00.7, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b1,     8'b11100001}, // D.01.7, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b1,     8'b11100010}, // D.02.7, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b0,     8'b11110011}, // D.19.7, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b1,     8'b11100100}, // D.04.7, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b0,     8'b11110101}, // D.21.7, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b0,     8'b11110110}, // D.22.7, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b1,     1'b0,     1'b1,     1'b1,     8'b11110111}, // K.23.7, disp_front = 1, disp_end = 1, K = 1, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b1,     8'b11101000}, // D.08.7, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b0,     8'b11111001}, // D.25.7, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b0,     8'b11111010}, // D.26.7, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b1,     1'b0,     1'b1,     1'b1,     8'b11111011}, // K.27.7, disp_front = 1, disp_end = 1, K = 1, code_err = 0, disp_err = 1
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b0,     8'b11111100}, // D.28.7, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b1,     1'b0,     1'b1,     1'b1,     8'b11111101}, // K.29.7, disp_front = 1, disp_end = 1, K = 1, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b0,     1'b1,     1'b1,     8'b11111110}, // K.30.7, disp_front = 1, disp_end = 1, K = 1, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b1,     8'b11100000}, // D.00.7, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b1,     8'b11100000}, // D.00.7, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b1,     8'b11111110}, // D.30.7, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b1,     8'b11111101}, // D.29.7, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b0,     8'b11100011}, // D.03.7, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b1,     8'b11111011}, // D.27.7, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b0,     8'b11100101}, // D.05.7, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b0,     8'b11100110}, // D.06.7, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b1,     8'b11101000}, // D.08.7, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b1,     8'b11110111}, // D.23.7, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b0,     8'b11101001}, // D.09.7, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b0,     8'b11101010}, // D.10.7, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b1,     8'b11100100}, // D.04.7, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b0,     8'b11101100}, // D.12.7, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b1,     8'b11100010}, // D.02.7, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b1,     8'b11100001}, // D.01.7, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b1,     8'b11100000}, // D.00.7, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b1,     8'b11100000}, // D.00.7, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b0,     8'b11110001}, // D.17.7, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b0,     8'b11110010}, // D.18.7, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b1,     8'b11111000}, // D.24.7, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b0,     8'b11110100}, // D.20.7, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b1,     8'b11111111}, // D.31.7, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b1,     8'b11110000}, // D.16.7, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b1,     8'b11100000}, // D.00.7, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b0,     8'b11100111}, // D.07.7, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b1,     8'b11100000}, // D.00.7, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b1,     8'b11101111}, // D.15.7, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b1,     8'b11100000}, // D.00.7, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b0,     1'b1,     1'b1,     8'b11111100}, // K.28.7, disp_front = 1, disp_end = 1, K = 1, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b1,     8'b11100000}, // D.00.7, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b1,     8'b11100000}, // D.00.7, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b1,     8'b11100000}, // D.00.7, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b1,     8'b00000000}, // D.00.0, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b1,     8'b00000000}, // D.00.0, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b1,     8'b00000000}, // D.00.0, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b1,     8'b00011100}, // D.28.0, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b1,     8'b00000000}, // D.00.0, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b1,     8'b00001111}, // D.15.0, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b1,     8'b00000000}, // D.00.0, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b0,     8'b00000111}, // D.07.0, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b1,     8'b00000000}, // D.00.0, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b1,     8'b00010000}, // D.16.0, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b1,     8'b00011111}, // D.31.0, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b0,     8'b00001011}, // D.11.0, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b1,     8'b00011000}, // D.24.0, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b0,     8'b00001101}, // D.13.0, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b0,     8'b00001110}, // D.14.0, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b1,     8'b00000000}, // D.00.0, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b1,     8'b00000000}, // D.00.0, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b1,     8'b00000001}, // D.01.0, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b1,     8'b00000010}, // D.02.0, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b0,     8'b00010011}, // D.19.0, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b1,     8'b00000100}, // D.04.0, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b0,     8'b00010101}, // D.21.0, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b0,     8'b00010110}, // D.22.0, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b1,     8'b00010111}, // D.23.0, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b1,     8'b00001000}, // D.08.0, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b0,     8'b00011001}, // D.25.0, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b0,     8'b00011010}, // D.26.0, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b1,     8'b00011011}, // D.27.0, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b0,     8'b00011100}, // D.28.0, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b1,     8'b00011101}, // D.29.0, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b1,     8'b00011110}, // D.30.0, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b1,     8'b00000000}, // D.00.0, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b1,     8'b00000000}, // D.00.0, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b1,     8'b00011110}, // D.30.0, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b1,     8'b00011101}, // D.29.0, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b0,     8'b00000011}, // D.03.0, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b1,     8'b00011011}, // D.27.0, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b0,     8'b00000101}, // D.05.0, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b0,     8'b00000110}, // D.06.0, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b1,     8'b00001000}, // D.08.0, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b1,     8'b00010111}, // D.23.0, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b0,     8'b00001001}, // D.09.0, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b0,     8'b00001010}, // D.10.0, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b1,     8'b00000100}, // D.04.0, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b0,     8'b00001100}, // D.12.0, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b1,     8'b00000010}, // D.02.0, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b1,     8'b00000001}, // D.01.0, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b1,     8'b00000000}, // D.00.0, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b1,     8'b00000000}, // D.00.0, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b0,     8'b00010001}, // D.17.0, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b0,     8'b00010010}, // D.18.0, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b1,     8'b00011000}, // D.24.0, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b0,     8'b00010100}, // D.20.0, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b1,     8'b00011111}, // D.31.0, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b1,     8'b00010000}, // D.16.0, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b1,     8'b00000000}, // D.00.0, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b0,     8'b00000111}, // D.07.0, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b1,     8'b00000000}, // D.00.0, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b1,     8'b00001111}, // D.15.0, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b1,     8'b00000000}, // D.00.0, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b0,     1'b1,     1'b1,     8'b00011100}, // K.28.0, disp_front = 1, disp_end = 1, K = 1, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b1,     8'b00000000}, // D.00.0, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b1,     8'b00000000}, // D.00.0, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b1,     8'b00000000}, // D.00.0, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b0,     8'b01100000}, // D.00.3, disp_front = 1, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b0,     8'b01100000}, // D.00.3, disp_front = 1, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b0,     8'b01100000}, // D.00.3, disp_front = 1, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b0,     1'b0,     1'b1,     1'b0,     8'b01111100}, // K.28.3, disp_front = 1, disp_end = 0, K = 1, code_err = 0, disp_err = 0
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b0,     8'b01100000}, // D.00.3, disp_front = 1, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b0,     8'b01101111}, // D.15.3, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b0,     8'b01100000}, // D.00.3, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b1,     8'b01100111}, // D.07.3, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b0,     8'b01100000}, // D.00.3, disp_front = 1, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b0,     8'b01110000}, // D.16.3, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b0,     8'b01111111}, // D.31.3, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b1,     8'b01101011}, // D.11.3, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b0,     8'b01111000}, // D.24.3, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b1,     8'b01101101}, // D.13.3, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b1,     8'b01101110}, // D.14.3, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b0,     8'b01100000}, // D.00.3, disp_front = 1, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b0,     8'b01100000}, // D.00.3, disp_front = 1, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b0,     8'b01100001}, // D.01.3, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b0,     8'b01100010}, // D.02.3, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b1,     8'b01110011}, // D.19.3, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b0,     8'b01100100}, // D.04.3, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b1,     8'b01110101}, // D.21.3, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b1,     8'b01110110}, // D.22.3, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b0,     8'b01110111}, // D.23.3, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b0,     8'b01101000}, // D.08.3, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b1,     8'b01111001}, // D.25.3, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b1,     8'b01111010}, // D.26.3, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b0,     8'b01111011}, // D.27.3, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b1,     8'b01111100}, // D.28.3, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b0,     8'b01111101}, // D.29.3, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b0,     8'b01111110}, // D.30.3, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b0,     8'b01100000}, // D.00.3, disp_front = 1, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b0,     8'b01100000}, // D.00.3, disp_front = 1, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b0,     8'b01111110}, // D.30.3, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b0,     8'b01111101}, // D.29.3, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b1,     8'b01100011}, // D.03.3, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b0,     8'b01111011}, // D.27.3, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b1,     8'b01100101}, // D.05.3, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b1,     8'b01100110}, // D.06.3, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b0,     8'b01101000}, // D.08.3, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b0,     8'b01110111}, // D.23.3, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b1,     8'b01101001}, // D.09.3, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b1,     8'b01101010}, // D.10.3, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b0,     8'b01100100}, // D.04.3, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b1,     8'b01101100}, // D.12.3, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b0,     8'b01100010}, // D.02.3, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b0,     8'b01100001}, // D.01.3, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b0,     8'b01100000}, // D.00.3, disp_front = 1, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b0,     1'b1,     1'b0,     1'b0,     8'b01100000}, // D.00.3, disp_front = 1, disp_end = 0, K = 0, code_err = 1, disp_err = 0
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b1,     8'b01110001}, // D.17.3, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b1,     8'b01110010}, // D.18.3, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b0,     8'b01111000}, // D.24.3, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b1,     8'b01110100}, // D.20.3, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b0,     8'b01111111}, // D.31.3, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b0,     8'b01110000}, // D.16.3, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b0,     8'b01100000}, // D.00.3, disp_front = 1, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b1,     8'b01100111}, // D.07.3, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b0,     8'b01100000}, // D.00.3, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b0,     8'b01101111}, // D.15.3, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b0,     8'b01100000}, // D.00.3, disp_front = 1, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b0,     8'b01111100}, // D.28.3, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b0,     8'b01100000}, // D.00.3, disp_front = 1, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b0,     8'b01100000}, // D.00.3, disp_front = 1, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b0,     8'b01100000}, // D.00.3, disp_front = 1, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b1,     8'b10000000}, // D.00.4, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b1,     8'b10000000}, // D.00.4, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b1,     8'b10000000}, // D.00.4, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b1,     8'b10011100}, // D.28.4, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b1,     8'b10000000}, // D.00.4, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b1,     8'b10001111}, // D.15.4, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b1,     8'b10000000}, // D.00.4, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b0,     8'b10000111}, // D.07.4, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b1,     8'b10000000}, // D.00.4, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b1,     8'b10010000}, // D.16.4, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b1,     8'b10011111}, // D.31.4, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b0,     8'b10001011}, // D.11.4, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b1,     8'b10011000}, // D.24.4, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b0,     8'b10001101}, // D.13.4, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b0,     8'b10001110}, // D.14.4, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b1,     8'b10000000}, // D.00.4, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b1,     8'b10000000}, // D.00.4, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b1,     8'b10000001}, // D.01.4, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b1,     8'b10000010}, // D.02.4, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b0,     8'b10010011}, // D.19.4, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b1,     8'b10000100}, // D.04.4, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b0,     8'b10010101}, // D.21.4, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b0,     8'b10010110}, // D.22.4, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b1,     8'b10010111}, // D.23.4, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b1,     8'b10001000}, // D.08.4, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b0,     8'b10011001}, // D.25.4, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b0,     8'b10011010}, // D.26.4, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b1,     8'b10011011}, // D.27.4, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b0,     8'b10011100}, // D.28.4, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b1,     8'b10011101}, // D.29.4, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b1,     8'b10011110}, // D.30.4, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b1,     8'b10000000}, // D.00.4, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b1,     8'b10000000}, // D.00.4, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b1,     8'b10011110}, // D.30.4, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b1,     8'b10011101}, // D.29.4, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b0,     8'b10000011}, // D.03.4, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b1,     8'b10011011}, // D.27.4, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b0,     8'b10000101}, // D.05.4, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b0,     8'b10000110}, // D.06.4, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b1,     8'b10001000}, // D.08.4, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b1,     8'b10010111}, // D.23.4, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b0,     8'b10001001}, // D.09.4, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b0,     8'b10001010}, // D.10.4, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b1,     8'b10000100}, // D.04.4, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b0,     8'b10001100}, // D.12.4, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b1,     8'b10000010}, // D.02.4, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b1,     8'b10000001}, // D.01.4, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b1,     8'b10000000}, // D.00.4, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b1,     8'b10000000}, // D.00.4, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b0,     8'b10010001}, // D.17.4, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b0,     8'b10010010}, // D.18.4, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b1,     8'b10011000}, // D.24.4, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b0,     8'b10010100}, // D.20.4, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b1,     8'b10011111}, // D.31.4, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b1,     8'b10010000}, // D.16.4, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b1,     8'b10000000}, // D.00.4, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b0,     8'b10000111}, // D.07.4, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b1,     8'b10000000}, // D.00.4, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b1,     8'b10001111}, // D.15.4, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b1,     8'b10000000}, // D.00.4, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b0,     1'b1,     1'b1,     8'b10011100}, // K.28.4, disp_front = 1, disp_end = 1, K = 1, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b1,     8'b10000000}, // D.00.4, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b1,     8'b10000000}, // D.00.4, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b1,     8'b10000000}, // D.00.4, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b0,     8'b10100000}, // D.00.5, disp_front = 1, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b0,     8'b10100000}, // D.00.5, disp_front = 1, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b0,     8'b10100000}, // D.00.5, disp_front = 1, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b0,     1'b0,     1'b1,     1'b0,     8'b01011100}, // K.28.2, disp_front = 1, disp_end = 0, K = 1, code_err = 0, disp_err = 0
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b0,     8'b10100000}, // D.00.5, disp_front = 1, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b0,     8'b10101111}, // D.15.5, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b0,     8'b10100000}, // D.00.5, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b1,     8'b10100111}, // D.07.5, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b0,     8'b10100000}, // D.00.5, disp_front = 1, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b0,     8'b10110000}, // D.16.5, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b0,     8'b10111111}, // D.31.5, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b1,     8'b10101011}, // D.11.5, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b0,     8'b10111000}, // D.24.5, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b1,     8'b10101101}, // D.13.5, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b1,     8'b10101110}, // D.14.5, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b0,     8'b10100000}, // D.00.5, disp_front = 1, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b0,     8'b10100000}, // D.00.5, disp_front = 1, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b0,     8'b10100001}, // D.01.5, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b0,     8'b10100010}, // D.02.5, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b1,     8'b10110011}, // D.19.5, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b0,     8'b10100100}, // D.04.5, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b1,     8'b10110101}, // D.21.5, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b1,     8'b10110110}, // D.22.5, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b0,     8'b10110111}, // D.23.5, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b0,     8'b10101000}, // D.08.5, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b1,     8'b10111001}, // D.25.5, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b1,     8'b10111010}, // D.26.5, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b0,     8'b10111011}, // D.27.5, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b1,     8'b10111100}, // D.28.5, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b0,     8'b10111101}, // D.29.5, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b0,     8'b10111110}, // D.30.5, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b0,     8'b10100000}, // D.00.5, disp_front = 1, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b0,     8'b10100000}, // D.00.5, disp_front = 1, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b0,     8'b10111110}, // D.30.5, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b0,     8'b10111101}, // D.29.5, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b1,     8'b10100011}, // D.03.5, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b0,     8'b10111011}, // D.27.5, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b1,     8'b10100101}, // D.05.5, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b1,     8'b10100110}, // D.06.5, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b0,     8'b10101000}, // D.08.5, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b0,     8'b10110111}, // D.23.5, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b1,     8'b10101001}, // D.09.5, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b1,     8'b10101010}, // D.10.5, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b0,     8'b10100100}, // D.04.5, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b1,     8'b10101100}, // D.12.5, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b0,     8'b10100010}, // D.02.5, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b0,     8'b10100001}, // D.01.5, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b0,     8'b10100000}, // D.00.5, disp_front = 1, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b0,     1'b1,     1'b0,     1'b0,     8'b10100000}, // D.00.5, disp_front = 1, disp_end = 0, K = 0, code_err = 1, disp_err = 0
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b1,     8'b10110001}, // D.17.5, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b1,     8'b10110010}, // D.18.5, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b0,     8'b10111000}, // D.24.5, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b1,     8'b10110100}, // D.20.5, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b0,     8'b10111111}, // D.31.5, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b0,     8'b10110000}, // D.16.5, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b0,     8'b10100000}, // D.00.5, disp_front = 1, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b1,     8'b10100111}, // D.07.5, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b0,     8'b10100000}, // D.00.5, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b0,     8'b10101111}, // D.15.5, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b0,     8'b10100000}, // D.00.5, disp_front = 1, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b0,     1'b1,     1'b0,     8'b01011100}, // K.28.2, disp_front = 1, disp_end = 0, K = 1, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b0,     8'b10100000}, // D.00.5, disp_front = 1, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b0,     8'b10100000}, // D.00.5, disp_front = 1, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b0,     8'b10100000}, // D.00.5, disp_front = 1, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b0,     8'b11000000}, // D.00.6, disp_front = 1, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b0,     8'b11000000}, // D.00.6, disp_front = 1, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b0,     8'b11000000}, // D.00.6, disp_front = 1, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b0,     1'b0,     1'b1,     1'b0,     8'b00111100}, // K.28.1, disp_front = 1, disp_end = 0, K = 1, code_err = 0, disp_err = 0
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b0,     8'b11000000}, // D.00.6, disp_front = 1, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b0,     8'b11001111}, // D.15.6, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b0,     8'b11000000}, // D.00.6, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b1,     8'b11000111}, // D.07.6, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b0,     8'b11000000}, // D.00.6, disp_front = 1, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b0,     8'b11010000}, // D.16.6, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b0,     8'b11011111}, // D.31.6, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b1,     8'b11001011}, // D.11.6, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b0,     8'b11011000}, // D.24.6, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b1,     8'b11001101}, // D.13.6, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b1,     8'b11001110}, // D.14.6, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b0,     8'b11000000}, // D.00.6, disp_front = 1, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b0,     8'b11000000}, // D.00.6, disp_front = 1, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b0,     8'b11000001}, // D.01.6, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b0,     8'b11000010}, // D.02.6, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b1,     8'b11010011}, // D.19.6, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b0,     8'b11000100}, // D.04.6, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b1,     8'b11010101}, // D.21.6, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b1,     8'b11010110}, // D.22.6, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b0,     8'b11010111}, // D.23.6, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b0,     8'b11001000}, // D.08.6, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b1,     8'b11011001}, // D.25.6, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b1,     8'b11011010}, // D.26.6, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b0,     8'b11011011}, // D.27.6, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b1,     8'b11011100}, // D.28.6, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b0,     8'b11011101}, // D.29.6, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b0,     8'b11011110}, // D.30.6, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b0,     8'b11000000}, // D.00.6, disp_front = 1, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b0,     8'b11000000}, // D.00.6, disp_front = 1, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b0,     8'b11011110}, // D.30.6, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b0,     8'b11011101}, // D.29.6, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b1,     8'b11000011}, // D.03.6, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b0,     8'b11011011}, // D.27.6, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b1,     8'b11000101}, // D.05.6, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b1,     8'b11000110}, // D.06.6, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b0,     8'b11001000}, // D.08.6, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b0,     8'b11010111}, // D.23.6, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b1,     8'b11001001}, // D.09.6, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b1,     8'b11001010}, // D.10.6, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b0,     8'b11000100}, // D.04.6, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b1,     8'b11001100}, // D.12.6, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b0,     8'b11000010}, // D.02.6, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b0,     8'b11000001}, // D.01.6, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b0,     8'b11000000}, // D.00.6, disp_front = 1, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b0,     1'b1,     1'b0,     1'b0,     8'b11000000}, // D.00.6, disp_front = 1, disp_end = 0, K = 0, code_err = 1, disp_err = 0
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b1,     8'b11010001}, // D.17.6, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b1,     8'b11010010}, // D.18.6, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b0,     8'b11011000}, // D.24.6, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b1,     8'b11010100}, // D.20.6, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b0,     8'b11011111}, // D.31.6, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b0,     8'b11010000}, // D.16.6, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b0,     8'b11000000}, // D.00.6, disp_front = 1, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b1,     8'b11000111}, // D.07.6, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b0,     8'b11000000}, // D.00.6, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b0,     8'b11001111}, // D.15.6, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b0,     8'b11000000}, // D.00.6, disp_front = 1, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b0,     1'b1,     1'b0,     8'b00111100}, // K.28.1, disp_front = 1, disp_end = 0, K = 1, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b0,     8'b11000000}, // D.00.6, disp_front = 1, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b0,     8'b11000000}, // D.00.6, disp_front = 1, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b0,     8'b11000000}, // D.00.6, disp_front = 1, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b1,     8'b11100000}, // D.00.7, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b1,     8'b11100000}, // D.00.7, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b1,     8'b11100000}, // D.00.7, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b1,     8'b11111100}, // D.28.7, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b1,     8'b11100000}, // D.00.7, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b1,     8'b11101111}, // D.15.7, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b1,     8'b11100000}, // D.00.7, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b0,     8'b11100111}, // D.07.7, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b1,     8'b11100000}, // D.00.7, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b1,     8'b11110000}, // D.16.7, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b1,     8'b11111111}, // D.31.7, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b0,     8'b11101011}, // D.11.7, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b1,     8'b11111000}, // D.24.7, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b0,     8'b11101101}, // D.13.7, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b0,     8'b11101110}, // D.14.7, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b1,     8'b11100000}, // D.00.7, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b1,     8'b11100000}, // D.00.7, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b1,     8'b11100001}, // D.01.7, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b1,     8'b11100010}, // D.02.7, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b0,     8'b11110011}, // D.19.7, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b1,     8'b11100100}, // D.04.7, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b0,     8'b11110101}, // D.21.7, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b0,     8'b11110110}, // D.22.7, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b1,     8'b11110111}, // D.23.7, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b1,     8'b11101000}, // D.08.7, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b0,     8'b11111001}, // D.25.7, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b0,     8'b11111010}, // D.26.7, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b1,     8'b11111011}, // D.27.7, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b0,     8'b11111100}, // D.28.7, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b1,     8'b11111101}, // D.29.7, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b1,     8'b11111110}, // D.30.7, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b1,     8'b11100000}, // D.00.7, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b1,     8'b11100000}, // D.00.7, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b1,     8'b11111110}, // D.30.7, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b1,     8'b11111101}, // D.29.7, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b0,     8'b11100011}, // D.03.7, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b1,     8'b11111011}, // D.27.7, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b0,     8'b11100101}, // D.05.7, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b0,     8'b11100110}, // D.06.7, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b1,     8'b11101000}, // D.08.7, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b1,     8'b11110111}, // D.23.7, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b0,     8'b11101001}, // D.09.7, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b0,     8'b11101010}, // D.10.7, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b1,     8'b11100100}, // D.04.7, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b0,     8'b11101100}, // D.12.7, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b1,     8'b11100010}, // D.02.7, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b1,     8'b11100001}, // D.01.7, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b1,     8'b11100000}, // D.00.7, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b0,     1'b1,     1'b0,     1'b1,     8'b11100000}, // D.00.7, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 0
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b0,     8'b11110001}, // D.17.7, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b0,     8'b11110010}, // D.18.7, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b1,     8'b11111000}, // D.24.7, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b0,     8'b11110100}, // D.20.7, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b1,     8'b11111111}, // D.31.7, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b1,     8'b11110000}, // D.16.7, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b1,     8'b11100000}, // D.00.7, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b0,     8'b11100111}, // D.07.7, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b1,     8'b11100000}, // D.00.7, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b1,     8'b11101111}, // D.15.7, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b1,     8'b11100000}, // D.00.7, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b1,     8'b11111100}, // D.28.7, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b1,     8'b11100000}, // D.00.7, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b1,     8'b11100000}, // D.00.7, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b1,     8'b11100000}, // D.00.7, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b1,     8'b11100000}, // D.00.7, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b1,     8'b11100000}, // D.00.7, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b1,     8'b11100000}, // D.00.7, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b1,     8'b11111100}, // D.28.7, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b1,     8'b11100000}, // D.00.7, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b1,     8'b11101111}, // D.15.7, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b1,     8'b11100000}, // D.00.7, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b0,     8'b11100111}, // D.07.7, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b1,     8'b11100000}, // D.00.7, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b1,     8'b11110000}, // D.16.7, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b1,     8'b11111111}, // D.31.7, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b0,     8'b11101011}, // D.11.7, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b1,     8'b11111000}, // D.24.7, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b0,     8'b11101101}, // D.13.7, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b0,     8'b11101110}, // D.14.7, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b1,     8'b11100000}, // D.00.7, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b1,     8'b11100000}, // D.00.7, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b1,     8'b11100001}, // D.01.7, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b1,     8'b11100010}, // D.02.7, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b0,     8'b11110011}, // D.19.7, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b1,     8'b11100100}, // D.04.7, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b0,     8'b11110101}, // D.21.7, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b0,     8'b11110110}, // D.22.7, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b1,     8'b11110111}, // D.23.7, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b1,     8'b11101000}, // D.08.7, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b0,     8'b11111001}, // D.25.7, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b0,     8'b11111010}, // D.26.7, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b1,     8'b11111011}, // D.27.7, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b0,     8'b11111100}, // D.28.7, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b1,     8'b11111101}, // D.29.7, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b1,     8'b11111110}, // D.30.7, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b1,     8'b11100000}, // D.00.7, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b1,     8'b11100000}, // D.00.7, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b1,     8'b11111110}, // D.30.7, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b1,     8'b11111101}, // D.29.7, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b0,     8'b11100011}, // D.03.7, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b1,     8'b11111011}, // D.27.7, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b0,     8'b11100101}, // D.05.7, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b0,     8'b11100110}, // D.06.7, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b1,     8'b11101000}, // D.08.7, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b1,     8'b11110111}, // D.23.7, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b0,     8'b11101001}, // D.09.7, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b0,     8'b11101010}, // D.10.7, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b1,     8'b11100100}, // D.04.7, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b0,     8'b11101100}, // D.12.7, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b1,     8'b11100010}, // D.02.7, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b1,     8'b11100001}, // D.01.7, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b1,     8'b11100000}, // D.00.7, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b1,     8'b11100000}, // D.00.7, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b0,     8'b11110001}, // D.17.7, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b0,     8'b11110010}, // D.18.7, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b1,     8'b11111000}, // D.24.7, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b0,     8'b11110100}, // D.20.7, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b1,     8'b11111111}, // D.31.7, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b1,     8'b11110000}, // D.16.7, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b1,     8'b11100000}, // D.00.7, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b0,     8'b11100111}, // D.07.7, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b1,     8'b11100000}, // D.00.7, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b1,     8'b11101111}, // D.15.7, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b1,     8'b11100000}, // D.00.7, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b1,     8'b11111100}, // D.28.7, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b1,     8'b11100000}, // D.00.7, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b1,     8'b11100000}, // D.00.7, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b1,     8'b11100000}, // D.00.7, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b0,     8'b00100000}, // D.00.1, disp_front = 1, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b0,     8'b00100000}, // D.00.1, disp_front = 1, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b0,     8'b00100000}, // D.00.1, disp_front = 1, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b0,     1'b0,     1'b1,     1'b0,     8'b11011100}, // K.28.6, disp_front = 1, disp_end = 0, K = 1, code_err = 0, disp_err = 0
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b0,     8'b00100000}, // D.00.1, disp_front = 1, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b0,     8'b00101111}, // D.15.1, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b0,     8'b00100000}, // D.00.1, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b1,     8'b00100111}, // D.07.1, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b0,     8'b00100000}, // D.00.1, disp_front = 1, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b0,     8'b00110000}, // D.16.1, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b0,     8'b00111111}, // D.31.1, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b1,     8'b00101011}, // D.11.1, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b0,     8'b00111000}, // D.24.1, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b1,     8'b00101101}, // D.13.1, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b1,     8'b00101110}, // D.14.1, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b0,     8'b00100000}, // D.00.1, disp_front = 1, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b0,     8'b00100000}, // D.00.1, disp_front = 1, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b0,     8'b00100001}, // D.01.1, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b0,     8'b00100010}, // D.02.1, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b1,     8'b00110011}, // D.19.1, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b0,     8'b00100100}, // D.04.1, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b1,     8'b00110101}, // D.21.1, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b1,     8'b00110110}, // D.22.1, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b0,     8'b00110111}, // D.23.1, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b0,     8'b00101000}, // D.08.1, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b1,     8'b00111001}, // D.25.1, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b1,     8'b00111010}, // D.26.1, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b0,     8'b00111011}, // D.27.1, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b1,     8'b00111100}, // D.28.1, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b0,     8'b00111101}, // D.29.1, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b0,     8'b00111110}, // D.30.1, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b0,     8'b00100000}, // D.00.1, disp_front = 1, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b0,     8'b00100000}, // D.00.1, disp_front = 1, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b0,     8'b00111110}, // D.30.1, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b0,     8'b00111101}, // D.29.1, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b1,     8'b00100011}, // D.03.1, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b0,     8'b00111011}, // D.27.1, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b1,     8'b00100101}, // D.05.1, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b1,     8'b00100110}, // D.06.1, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b0,     8'b00101000}, // D.08.1, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b0,     8'b00110111}, // D.23.1, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b1,     8'b00101001}, // D.09.1, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b1,     8'b00101010}, // D.10.1, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b0,     8'b00100100}, // D.04.1, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b1,     8'b00101100}, // D.12.1, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b0,     8'b00100010}, // D.02.1, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b0,     8'b00100001}, // D.01.1, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b0,     8'b00100000}, // D.00.1, disp_front = 1, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b0,     1'b1,     1'b0,     1'b0,     8'b00100000}, // D.00.1, disp_front = 1, disp_end = 0, K = 0, code_err = 1, disp_err = 0
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b1,     8'b00110001}, // D.17.1, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b1,     8'b00110010}, // D.18.1, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b0,     8'b00111000}, // D.24.1, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b1,     8'b00110100}, // D.20.1, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b0,     8'b00111111}, // D.31.1, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b0,     8'b00110000}, // D.16.1, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b0,     8'b00100000}, // D.00.1, disp_front = 1, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b1,     8'b00100111}, // D.07.1, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b0,     8'b00100000}, // D.00.1, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b0,     8'b00101111}, // D.15.1, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b0,     8'b00100000}, // D.00.1, disp_front = 1, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b0,     1'b1,     1'b0,     8'b11011100}, // K.28.6, disp_front = 1, disp_end = 0, K = 1, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b0,     8'b00100000}, // D.00.1, disp_front = 1, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b0,     8'b00100000}, // D.00.1, disp_front = 1, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b0,     8'b00100000}, // D.00.1, disp_front = 1, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b0,     8'b01000000}, // D.00.2, disp_front = 1, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b0,     8'b01000000}, // D.00.2, disp_front = 1, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b0,     8'b01000000}, // D.00.2, disp_front = 1, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b0,     1'b0,     1'b1,     1'b0,     8'b10111100}, // K.28.5, disp_front = 1, disp_end = 0, K = 1, code_err = 0, disp_err = 0
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b0,     8'b01000000}, // D.00.2, disp_front = 1, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b0,     8'b01001111}, // D.15.2, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b0,     8'b01000000}, // D.00.2, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b1,     8'b01000111}, // D.07.2, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b0,     8'b01000000}, // D.00.2, disp_front = 1, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b0,     8'b01010000}, // D.16.2, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b0,     8'b01011111}, // D.31.2, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b1,     8'b01001011}, // D.11.2, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b0,     8'b01011000}, // D.24.2, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b1,     8'b01001101}, // D.13.2, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b1,     8'b01001110}, // D.14.2, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b0,     8'b01000000}, // D.00.2, disp_front = 1, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b0,     8'b01000000}, // D.00.2, disp_front = 1, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b0,     8'b01000001}, // D.01.2, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b0,     8'b01000010}, // D.02.2, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b1,     8'b01010011}, // D.19.2, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b0,     8'b01000100}, // D.04.2, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b1,     8'b01010101}, // D.21.2, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b1,     8'b01010110}, // D.22.2, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b0,     8'b01010111}, // D.23.2, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b0,     8'b01001000}, // D.08.2, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b1,     8'b01011001}, // D.25.2, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b1,     8'b01011010}, // D.26.2, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b0,     8'b01011011}, // D.27.2, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b1,     8'b01011100}, // D.28.2, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b0,     8'b01011101}, // D.29.2, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b0,     8'b01011110}, // D.30.2, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b0,     8'b01000000}, // D.00.2, disp_front = 1, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b0,     8'b01000000}, // D.00.2, disp_front = 1, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b0,     8'b01011110}, // D.30.2, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b0,     8'b01011101}, // D.29.2, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b1,     8'b01000011}, // D.03.2, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b0,     8'b01011011}, // D.27.2, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b1,     8'b01000101}, // D.05.2, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b1,     8'b01000110}, // D.06.2, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b0,     8'b01001000}, // D.08.2, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b0,     8'b01010111}, // D.23.2, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b1,     8'b01001001}, // D.09.2, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b1,     8'b01001010}, // D.10.2, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b0,     8'b01000100}, // D.04.2, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b1,     8'b01001100}, // D.12.2, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b0,     8'b01000010}, // D.02.2, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b0,     8'b01000001}, // D.01.2, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b0,     8'b01000000}, // D.00.2, disp_front = 1, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b0,     1'b1,     1'b0,     1'b0,     8'b01000000}, // D.00.2, disp_front = 1, disp_end = 0, K = 0, code_err = 1, disp_err = 0
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b1,     8'b01010001}, // D.17.2, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b1,     8'b01010010}, // D.18.2, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b0,     8'b01011000}, // D.24.2, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b1,     8'b01010100}, // D.20.2, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b0,     8'b01011111}, // D.31.2, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b0,     8'b01010000}, // D.16.2, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b0,     8'b01000000}, // D.00.2, disp_front = 1, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b1,     8'b01000111}, // D.07.2, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b0,     8'b01000000}, // D.00.2, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b0,     8'b01001111}, // D.15.2, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b0,     8'b01000000}, // D.00.2, disp_front = 1, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b0,     1'b1,     1'b0,     8'b10111100}, // K.28.5, disp_front = 1, disp_end = 0, K = 1, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b0,     8'b01000000}, // D.00.2, disp_front = 1, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b0,     8'b01000000}, // D.00.2, disp_front = 1, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b0,     8'b01000000}, // D.00.2, disp_front = 1, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b1,     8'b10000000}, // D.00.4, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b1,     8'b10000000}, // D.00.4, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b1,     8'b10000000}, // D.00.4, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b0,     1'b0,     1'b1,     1'b1,     8'b10011100}, // K.28.4, disp_front = 1, disp_end = 1, K = 1, code_err = 0, disp_err = 0
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b1,     8'b10000000}, // D.00.4, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b1,     8'b10001111}, // D.15.4, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b1,     8'b10000000}, // D.00.4, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b0,     8'b10000111}, // D.07.4, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b1,     8'b10000000}, // D.00.4, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b1,     8'b10010000}, // D.16.4, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b1,     8'b10011111}, // D.31.4, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b0,     8'b10001011}, // D.11.4, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b1,     8'b10011000}, // D.24.4, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b0,     8'b10001101}, // D.13.4, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b0,     8'b10001110}, // D.14.4, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b1,     8'b10000000}, // D.00.4, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b1,     8'b10000000}, // D.00.4, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b1,     8'b10000001}, // D.01.4, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b1,     8'b10000010}, // D.02.4, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b0,     8'b10010011}, // D.19.4, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b1,     8'b10000100}, // D.04.4, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b0,     8'b10010101}, // D.21.4, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b0,     8'b10010110}, // D.22.4, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b1,     8'b10010111}, // D.23.4, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b1,     8'b10001000}, // D.08.4, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b0,     8'b10011001}, // D.25.4, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b0,     8'b10011010}, // D.26.4, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b1,     8'b10011011}, // D.27.4, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b0,     8'b10011100}, // D.28.4, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b1,     8'b10011101}, // D.29.4, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b1,     8'b10011110}, // D.30.4, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b1,     8'b10000000}, // D.00.4, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b1,     8'b10000000}, // D.00.4, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b1,     8'b10011110}, // D.30.4, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b1,     8'b10011101}, // D.29.4, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b0,     8'b10000011}, // D.03.4, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b1,     8'b10011011}, // D.27.4, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b0,     8'b10000101}, // D.05.4, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b0,     8'b10000110}, // D.06.4, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b1,     8'b10001000}, // D.08.4, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b1,     8'b10010111}, // D.23.4, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b0,     8'b10001001}, // D.09.4, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b0,     8'b10001010}, // D.10.4, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b1,     8'b10000100}, // D.04.4, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b0,     8'b10001100}, // D.12.4, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b1,     8'b10000010}, // D.02.4, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b1,     8'b10000001}, // D.01.4, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b1,     8'b10000000}, // D.00.4, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b0,     1'b1,     1'b0,     1'b1,     8'b10000000}, // D.00.4, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 0
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b0,     8'b10010001}, // D.17.4, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b0,     8'b10010010}, // D.18.4, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b1,     8'b10011000}, // D.24.4, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b0,     8'b10010100}, // D.20.4, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b1,     8'b10011111}, // D.31.4, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b1,     8'b10010000}, // D.16.4, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b1,     8'b10000000}, // D.00.4, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b0,     8'b10000111}, // D.07.4, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b1,     8'b10000000}, // D.00.4, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b1,     8'b10001111}, // D.15.4, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b1,     8'b10000000}, // D.00.4, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b1,     8'b10011100}, // D.28.4, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b1,     8'b10000000}, // D.00.4, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b1,     8'b10000000}, // D.00.4, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b1,     8'b10000000}, // D.00.4, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b0,     8'b01100000}, // D.00.3, disp_front = 1, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b0,     8'b01100000}, // D.00.3, disp_front = 1, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b0,     8'b01100000}, // D.00.3, disp_front = 1, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b0,     8'b01111100}, // D.28.3, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b0,     8'b01100000}, // D.00.3, disp_front = 1, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b0,     8'b01101111}, // D.15.3, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b0,     8'b01100000}, // D.00.3, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b1,     8'b01100111}, // D.07.3, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b0,     8'b01100000}, // D.00.3, disp_front = 1, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b0,     8'b01110000}, // D.16.3, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b0,     8'b01111111}, // D.31.3, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b1,     8'b01101011}, // D.11.3, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b0,     8'b01111000}, // D.24.3, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b1,     8'b01101101}, // D.13.3, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b1,     8'b01101110}, // D.14.3, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b0,     8'b01100000}, // D.00.3, disp_front = 1, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b0,     8'b01100000}, // D.00.3, disp_front = 1, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b0,     8'b01100001}, // D.01.3, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b0,     8'b01100010}, // D.02.3, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b1,     8'b01110011}, // D.19.3, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b0,     8'b01100100}, // D.04.3, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b1,     8'b01110101}, // D.21.3, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b1,     8'b01110110}, // D.22.3, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b0,     8'b01110111}, // D.23.3, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b0,     8'b01101000}, // D.08.3, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b1,     8'b01111001}, // D.25.3, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b1,     8'b01111010}, // D.26.3, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b0,     8'b01111011}, // D.27.3, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b1,     8'b01111100}, // D.28.3, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b0,     8'b01111101}, // D.29.3, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b0,     8'b01111110}, // D.30.3, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b0,     8'b01100000}, // D.00.3, disp_front = 1, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b0,     8'b01100000}, // D.00.3, disp_front = 1, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b0,     8'b01111110}, // D.30.3, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b0,     8'b01111101}, // D.29.3, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b1,     8'b01100011}, // D.03.3, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b0,     8'b01111011}, // D.27.3, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b1,     8'b01100101}, // D.05.3, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b1,     8'b01100110}, // D.06.3, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b0,     8'b01101000}, // D.08.3, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b0,     8'b01110111}, // D.23.3, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b1,     8'b01101001}, // D.09.3, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b1,     8'b01101010}, // D.10.3, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b0,     8'b01100100}, // D.04.3, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b1,     8'b01101100}, // D.12.3, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b0,     8'b01100010}, // D.02.3, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b0,     8'b01100001}, // D.01.3, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b0,     8'b01100000}, // D.00.3, disp_front = 1, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b0,     1'b1,     1'b0,     1'b0,     8'b01100000}, // D.00.3, disp_front = 1, disp_end = 0, K = 0, code_err = 1, disp_err = 0
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b1,     8'b01110001}, // D.17.3, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b1,     8'b01110010}, // D.18.3, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b0,     8'b01111000}, // D.24.3, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b1,     8'b01110100}, // D.20.3, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b0,     8'b01111111}, // D.31.3, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b0,     8'b01110000}, // D.16.3, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b0,     8'b01100000}, // D.00.3, disp_front = 1, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b1,     8'b01100111}, // D.07.3, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b0,     8'b01100000}, // D.00.3, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b0,     8'b01101111}, // D.15.3, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b0,     8'b01100000}, // D.00.3, disp_front = 1, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b0,     1'b1,     1'b0,     8'b01111100}, // K.28.3, disp_front = 1, disp_end = 0, K = 1, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b0,     8'b01100000}, // D.00.3, disp_front = 1, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b0,     8'b01100000}, // D.00.3, disp_front = 1, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b0,     8'b01100000}, // D.00.3, disp_front = 1, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b1,     8'b00000000}, // D.00.0, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b1,     8'b00000000}, // D.00.0, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b1,     8'b00000000}, // D.00.0, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b0,     1'b0,     1'b1,     1'b1,     8'b00011100}, // K.28.0, disp_front = 1, disp_end = 1, K = 1, code_err = 0, disp_err = 0
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b1,     8'b00000000}, // D.00.0, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b1,     8'b00001111}, // D.15.0, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b1,     8'b00000000}, // D.00.0, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b0,     8'b00000111}, // D.07.0, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b1,     8'b00000000}, // D.00.0, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b1,     8'b00010000}, // D.16.0, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b1,     8'b00011111}, // D.31.0, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b0,     8'b00001011}, // D.11.0, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b1,     8'b00011000}, // D.24.0, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b0,     8'b00001101}, // D.13.0, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b0,     8'b00001110}, // D.14.0, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b1,     8'b00000000}, // D.00.0, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b1,     8'b00000000}, // D.00.0, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b1,     8'b00000001}, // D.01.0, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b1,     8'b00000010}, // D.02.0, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b0,     8'b00010011}, // D.19.0, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b1,     8'b00000100}, // D.04.0, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b0,     8'b00010101}, // D.21.0, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b0,     8'b00010110}, // D.22.0, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b1,     8'b00010111}, // D.23.0, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b1,     8'b00001000}, // D.08.0, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b0,     8'b00011001}, // D.25.0, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b0,     8'b00011010}, // D.26.0, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b1,     8'b00011011}, // D.27.0, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b0,     8'b00011100}, // D.28.0, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b1,     8'b00011101}, // D.29.0, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b1,     8'b00011110}, // D.30.0, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b1,     8'b00000000}, // D.00.0, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b1,     8'b00000000}, // D.00.0, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b1,     8'b00011110}, // D.30.0, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b1,     8'b00011101}, // D.29.0, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b0,     8'b00000011}, // D.03.0, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b1,     8'b00011011}, // D.27.0, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b0,     8'b00000101}, // D.05.0, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b0,     8'b00000110}, // D.06.0, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b1,     8'b00001000}, // D.08.0, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b1,     8'b00010111}, // D.23.0, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b0,     8'b00001001}, // D.09.0, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b0,     8'b00001010}, // D.10.0, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b1,     8'b00000100}, // D.04.0, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b0,     8'b00001100}, // D.12.0, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b1,     8'b00000010}, // D.02.0, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b1,     8'b00000001}, // D.01.0, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b1,     8'b00000000}, // D.00.0, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b0,     1'b1,     1'b0,     1'b1,     8'b00000000}, // D.00.0, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 0
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b0,     8'b00010001}, // D.17.0, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b0,     8'b00010010}, // D.18.0, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b1,     8'b00011000}, // D.24.0, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b0,     8'b00010100}, // D.20.0, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b1,     8'b00011111}, // D.31.0, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b1,     8'b00010000}, // D.16.0, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b1,     8'b00000000}, // D.00.0, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b0,     8'b00000111}, // D.07.0, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b1,     8'b00000000}, // D.00.0, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b1,     8'b00001111}, // D.15.0, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b1,     8'b00000000}, // D.00.0, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b1,     8'b00011100}, // D.28.0, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b1,     8'b00000000}, // D.00.0, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b1,     8'b00000000}, // D.00.0, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b1,     8'b00000000}, // D.00.0, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b1,     8'b11100000}, // D.00.7, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b1,     8'b11100000}, // D.00.7, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b1,     8'b11100000}, // D.00.7, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b0,     1'b0,     1'b1,     1'b1,     8'b11111100}, // K.28.7, disp_front = 1, disp_end = 1, K = 1, code_err = 0, disp_err = 0
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b1,     8'b11100000}, // D.00.7, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b1,     8'b11101111}, // D.15.7, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b1,     8'b11100000}, // D.00.7, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b0,     8'b11100111}, // D.07.7, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b1,     8'b11100000}, // D.00.7, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b1,     8'b11110000}, // D.16.7, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b1,     8'b11111111}, // D.31.7, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b0,     8'b11101011}, // D.11.7, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b1,     8'b11111000}, // D.24.7, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b0,     8'b11101101}, // D.13.7, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b0,     8'b11101110}, // D.14.7, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b1,     8'b11100000}, // D.00.7, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b1,     8'b11100000}, // D.00.7, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b1,     8'b11100001}, // D.01.7, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b1,     8'b11100010}, // D.02.7, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b0,     8'b11110011}, // D.19.7, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b1,     8'b11100100}, // D.04.7, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b0,     8'b11110101}, // D.21.7, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b0,     8'b11110110}, // D.22.7, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b1,     8'b11110111}, // D.23.7, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b0,     1'b0,     1'b0,     1'b1,     8'b11101000}, // D.08.7, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 0
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b0,     8'b11111001}, // D.25.7, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b0,     8'b11111010}, // D.26.7, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b1,     8'b11111011}, // D.27.7, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b0,     8'b11111100}, // D.28.7, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b1,     8'b11111101}, // D.29.7, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b1,     8'b11111110}, // D.30.7, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b1,     8'b11100000}, // D.00.7, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b1,     8'b11100000}, // D.00.7, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b0,     1'b0,     1'b1,     1'b1,     8'b11111110}, // K.30.7, disp_front = 1, disp_end = 1, K = 1, code_err = 0, disp_err = 0
     {1'b1,       1'b0,     1'b0,     1'b1,     1'b1,     8'b11111101}, // K.29.7, disp_front = 1, disp_end = 1, K = 1, code_err = 0, disp_err = 0
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b0,     8'b11100011}, // D.03.7, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b0,     1'b0,     1'b1,     1'b1,     8'b11111011}, // K.27.7, disp_front = 1, disp_end = 1, K = 1, code_err = 0, disp_err = 0
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b0,     8'b11100101}, // D.05.7, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b0,     8'b11100110}, // D.06.7, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b1,     8'b11101000}, // D.08.7, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b0,     1'b0,     1'b1,     1'b1,     8'b11110111}, // K.23.7, disp_front = 1, disp_end = 1, K = 1, code_err = 0, disp_err = 0
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b0,     8'b11101001}, // D.09.7, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b0,     8'b11101010}, // D.10.7, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b1,     8'b11100100}, // D.04.7, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b0,     8'b11101100}, // D.12.7, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b1,     8'b11100010}, // D.02.7, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b1,     8'b11100001}, // D.01.7, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b1,     8'b11100000}, // D.00.7, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b0,     1'b1,     1'b0,     1'b1,     8'b11100000}, // D.00.7, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 0
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b0,     8'b11110001}, // D.17.7, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b0,     8'b11110010}, // D.18.7, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b1,     8'b11111000}, // D.24.7, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b0,     8'b11110100}, // D.20.7, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b1,     8'b11111111}, // D.31.7, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b1,     8'b11110000}, // D.16.7, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b1,     8'b11100000}, // D.00.7, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b0,     8'b11100111}, // D.07.7, disp_front = 1, disp_end = 0, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b1,     8'b11100000}, // D.00.7, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b1,     8'b11101111}, // D.15.7, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b1,     8'b11100000}, // D.00.7, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b0,     1'b0,     1'b1,     8'b11111100}, // D.28.7, disp_front = 1, disp_end = 1, K = 0, code_err = 0, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b1,     8'b11100000}, // D.00.7, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b1,     8'b11100000}, // D.00.7, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b1,     8'b11100000}, // D.00.7, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b1,     8'b00000000}, // D.00.0, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b1,     8'b00000000}, // D.00.0, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b1,     8'b00000000}, // D.00.0, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b1,     8'b00011100}, // D.28.0, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b1,     8'b00000000}, // D.00.0, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b1,     8'b00001111}, // D.15.0, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b1,     8'b00000000}, // D.00.0, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b0,     8'b00000111}, // D.07.0, disp_front = 1, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b1,     8'b00000000}, // D.00.0, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b1,     8'b00010000}, // D.16.0, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b1,     8'b00011111}, // D.31.0, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b0,     8'b00001011}, // D.11.0, disp_front = 1, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b1,     8'b00011000}, // D.24.0, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b0,     8'b00001101}, // D.13.0, disp_front = 1, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b0,     8'b00001110}, // D.14.0, disp_front = 1, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b1,     8'b00000000}, // D.00.0, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b1,     8'b00000000}, // D.00.0, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b1,     8'b00000001}, // D.01.0, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b1,     8'b00000010}, // D.02.0, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b0,     8'b00010011}, // D.19.0, disp_front = 1, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b1,     8'b00000100}, // D.04.0, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b0,     8'b00010101}, // D.21.0, disp_front = 1, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b0,     8'b00010110}, // D.22.0, disp_front = 1, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b1,     8'b00010111}, // D.23.0, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b1,     8'b00001000}, // D.08.0, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b0,     8'b00011001}, // D.25.0, disp_front = 1, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b0,     8'b00011010}, // D.26.0, disp_front = 1, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b1,     8'b00011011}, // D.27.0, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b0,     8'b00011100}, // D.28.0, disp_front = 1, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b1,     8'b00011101}, // D.29.0, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b1,     8'b00011110}, // D.30.0, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b1,     8'b00000000}, // D.00.0, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b1,     8'b00000000}, // D.00.0, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b1,     8'b00011110}, // D.30.0, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b1,     8'b00011101}, // D.29.0, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b0,     8'b00000011}, // D.03.0, disp_front = 1, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b1,     8'b00011011}, // D.27.0, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b0,     8'b00000101}, // D.05.0, disp_front = 1, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b0,     8'b00000110}, // D.06.0, disp_front = 1, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b1,     8'b00001000}, // D.08.0, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b1,     8'b00010111}, // D.23.0, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b0,     8'b00001001}, // D.09.0, disp_front = 1, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b0,     8'b00001010}, // D.10.0, disp_front = 1, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b1,     8'b00000100}, // D.04.0, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b0,     8'b00001100}, // D.12.0, disp_front = 1, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b1,     8'b00000010}, // D.02.0, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b1,     8'b00000001}, // D.01.0, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b1,     8'b00000000}, // D.00.0, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b1,     8'b00000000}, // D.00.0, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b0,     8'b00010001}, // D.17.0, disp_front = 1, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b0,     8'b00010010}, // D.18.0, disp_front = 1, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b1,     8'b00011000}, // D.24.0, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b0,     8'b00010100}, // D.20.0, disp_front = 1, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b1,     8'b00011111}, // D.31.0, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b1,     8'b00010000}, // D.16.0, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b1,     8'b00000000}, // D.00.0, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b0,     8'b00000111}, // D.07.0, disp_front = 1, disp_end = 0, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b1,     8'b00000000}, // D.00.0, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b1,     8'b00001111}, // D.15.0, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b1,     8'b00000000}, // D.00.0, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b1,     8'b00011100}, // D.28.0, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b1,     8'b00000000}, // D.00.0, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b1,     8'b00000000}, // D.00.0, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 1
     {1'b1,       1'b1,     1'b1,     1'b0,     1'b1,     8'b00000000}  // D.00.0, disp_front = 1, disp_end = 1, K = 0, code_err = 1, disp_err = 1
  };

endpackage