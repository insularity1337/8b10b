package pkg_8b10b;

  logic [1+1+2+8+10+2-1:0] enc_table [1024] = '{
  //WRONG K     RDF    octet        code            RDE
  //23    22    21:20  19:12        11:2            1:0
   {1'b0, 1'b0, 2'b11, 8'b00000000, 10'b1001110100, 2'b11}, // D00.0 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b00000000, 10'b0110001011, 2'b01}, // D00.0 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b00000001, 10'b0111010100, 2'b11}, // D01.0 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b00000001, 10'b1000101011, 2'b01}, // D01.0 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b00000010, 10'b1011010100, 2'b11}, // D02.0 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b00000010, 10'b0100101011, 2'b01}, // D02.0 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b00000011, 10'b1100011011, 2'b01}, // D03.0 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b00000011, 10'b1100010100, 2'b11}, // D03.0 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b00000100, 10'b1101010100, 2'b11}, // D04.0 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b00000100, 10'b0010101011, 2'b01}, // D04.0 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b00000101, 10'b1010011011, 2'b01}, // D05.0 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b00000101, 10'b1010010100, 2'b11}, // D05.0 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b00000110, 10'b0110011011, 2'b01}, // D06.0 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b00000110, 10'b0110010100, 2'b11}, // D06.0 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b00000111, 10'b1110001011, 2'b01}, // D07.0 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b00000111, 10'b0001110100, 2'b11}, // D07.0 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b00001000, 10'b1110010100, 2'b11}, // D08.0 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b00001000, 10'b0001101011, 2'b01}, // D08.0 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b00001001, 10'b1001011011, 2'b01}, // D09.0 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b00001001, 10'b1001010100, 2'b11}, // D09.0 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b00001010, 10'b0101011011, 2'b01}, // D10.0 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b00001010, 10'b0101010100, 2'b11}, // D10.0 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b00001011, 10'b1101001011, 2'b01}, // D11.0 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b00001011, 10'b1101000100, 2'b11}, // D11.0 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b00001100, 10'b0011011011, 2'b01}, // D12.0 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b00001100, 10'b0011010100, 2'b11}, // D12.0 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b00001101, 10'b1011001011, 2'b01}, // D13.0 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b00001101, 10'b1011000100, 2'b11}, // D13.0 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b00001110, 10'b0111001011, 2'b01}, // D14.0 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b00001110, 10'b0111000100, 2'b11}, // D14.0 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b00001111, 10'b0101110100, 2'b11}, // D15.0 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b00001111, 10'b1010001011, 2'b01}, // D15.0 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b00010000, 10'b0110110100, 2'b11}, // D16.0 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b00010000, 10'b1001001011, 2'b01}, // D16.0 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b00010001, 10'b1000111011, 2'b01}, // D17.0 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b00010001, 10'b1000110100, 2'b11}, // D17.0 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b00010010, 10'b0100111011, 2'b01}, // D18.0 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b00010010, 10'b0100110100, 2'b11}, // D18.0 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b00010011, 10'b1100101011, 2'b01}, // D19.0 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b00010011, 10'b1100100100, 2'b11}, // D19.0 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b00010100, 10'b0010111011, 2'b01}, // D20.0 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b00010100, 10'b0010110100, 2'b11}, // D20.0 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b00010101, 10'b1010101011, 2'b01}, // D21.0 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b00010101, 10'b1010100100, 2'b11}, // D21.0 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b00010110, 10'b0110101011, 2'b01}, // D22.0 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b00010110, 10'b0110100100, 2'b11}, // D22.0 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b00010111, 10'b1110100100, 2'b11}, // D23.0 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b00010111, 10'b0001011011, 2'b01}, // D23.0 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b00011000, 10'b1100110100, 2'b11}, // D24.0 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b00011000, 10'b0011001011, 2'b01}, // D24.0 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b00011001, 10'b1001101011, 2'b01}, // D25.0 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b00011001, 10'b1001100100, 2'b11}, // D25.0 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b00011010, 10'b0101101011, 2'b01}, // D26.0 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b00011010, 10'b0101100100, 2'b11}, // D26.0 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b00011011, 10'b1101100100, 2'b11}, // D27.0 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b00011011, 10'b0010011011, 2'b01}, // D27.0 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b00011100, 10'b0011101011, 2'b01}, // D28.0 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b00011100, 10'b0011100100, 2'b11}, // D28.0 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b00011101, 10'b1011100100, 2'b11}, // D29.0 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b00011101, 10'b0100011011, 2'b01}, // D29.0 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b00011110, 10'b0111100100, 2'b11}, // D30.0 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b00011110, 10'b1000011011, 2'b01}, // D30.0 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b00011111, 10'b1010110100, 2'b11}, // D31.0 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b00011111, 10'b0101001011, 2'b01}, // D31.0 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b00100000, 10'b1001111001, 2'b01}, // D00.1 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b00100000, 10'b0110001001, 2'b11}, // D00.1 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b00100001, 10'b0111011001, 2'b01}, // D01.1 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b00100001, 10'b1000101001, 2'b11}, // D01.1 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b00100010, 10'b1011011001, 2'b01}, // D02.1 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b00100010, 10'b0100101001, 2'b11}, // D02.1 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b00100011, 10'b1100011001, 2'b11}, // D03.1 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b00100011, 10'b1100011001, 2'b01}, // D03.1 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b00100100, 10'b1101011001, 2'b01}, // D04.1 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b00100100, 10'b0010101001, 2'b11}, // D04.1 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b00100101, 10'b1010011001, 2'b11}, // D05.1 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b00100101, 10'b1010011001, 2'b01}, // D05.1 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b00100110, 10'b0110011001, 2'b11}, // D06.1 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b00100110, 10'b0110011001, 2'b01}, // D06.1 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b00100111, 10'b1110001001, 2'b11}, // D07.1 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b00100111, 10'b0001111001, 2'b01}, // D07.1 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b00101000, 10'b1110011001, 2'b01}, // D08.1 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b00101000, 10'b0001101001, 2'b11}, // D08.1 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b00101001, 10'b1001011001, 2'b11}, // D09.1 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b00101001, 10'b1001011001, 2'b01}, // D09.1 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b00101010, 10'b0101011001, 2'b11}, // D10.1 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b00101010, 10'b0101011001, 2'b01}, // D10.1 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b00101011, 10'b1101001001, 2'b11}, // D11.1 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b00101011, 10'b1101001001, 2'b01}, // D11.1 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b00101100, 10'b0011011001, 2'b11}, // D12.1 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b00101100, 10'b0011011001, 2'b01}, // D12.1 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b00101101, 10'b1011001001, 2'b11}, // D13.1 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b00101101, 10'b1011001001, 2'b01}, // D13.1 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b00101110, 10'b0111001001, 2'b11}, // D14.1 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b00101110, 10'b0111001001, 2'b01}, // D14.1 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b00101111, 10'b0101111001, 2'b01}, // D15.1 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b00101111, 10'b1010001001, 2'b11}, // D15.1 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b00110000, 10'b0110111001, 2'b01}, // D16.1 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b00110000, 10'b1001001001, 2'b11}, // D16.1 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b00110001, 10'b1000111001, 2'b11}, // D17.1 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b00110001, 10'b1000111001, 2'b01}, // D17.1 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b00110010, 10'b0100111001, 2'b11}, // D18.1 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b00110010, 10'b0100111001, 2'b01}, // D18.1 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b00110011, 10'b1100101001, 2'b11}, // D19.1 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b00110011, 10'b1100101001, 2'b01}, // D19.1 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b00110100, 10'b0010111001, 2'b11}, // D20.1 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b00110100, 10'b0010111001, 2'b01}, // D20.1 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b00110101, 10'b1010101001, 2'b11}, // D21.1 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b00110101, 10'b1010101001, 2'b01}, // D21.1 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b00110110, 10'b0110101001, 2'b11}, // D22.1 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b00110110, 10'b0110101001, 2'b01}, // D22.1 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b00110111, 10'b1110101001, 2'b01}, // D23.1 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b00110111, 10'b0001011001, 2'b11}, // D23.1 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b00111000, 10'b1100111001, 2'b01}, // D24.1 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b00111000, 10'b0011001001, 2'b11}, // D24.1 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b00111001, 10'b1001101001, 2'b11}, // D25.1 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b00111001, 10'b1001101001, 2'b01}, // D25.1 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b00111010, 10'b0101101001, 2'b11}, // D26.1 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b00111010, 10'b0101101001, 2'b01}, // D26.1 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b00111011, 10'b1101101001, 2'b01}, // D27.1 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b00111011, 10'b0010011001, 2'b11}, // D27.1 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b00111100, 10'b0011101001, 2'b11}, // D28.1 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b00111100, 10'b0011101001, 2'b01}, // D28.1 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b00111101, 10'b1011101001, 2'b01}, // D29.1 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b00111101, 10'b0100011001, 2'b11}, // D29.1 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b00111110, 10'b0111101001, 2'b01}, // D30.1 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b00111110, 10'b1000011001, 2'b11}, // D30.1 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b00111111, 10'b1010111001, 2'b01}, // D31.1 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b00111111, 10'b0101001001, 2'b11}, // D31.1 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b01000000, 10'b1001110101, 2'b01}, // D00.2 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b01000000, 10'b0110000101, 2'b11}, // D00.2 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b01000001, 10'b0111010101, 2'b01}, // D01.2 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b01000001, 10'b1000100101, 2'b11}, // D01.2 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b01000010, 10'b1011010101, 2'b01}, // D02.2 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b01000010, 10'b0100100101, 2'b11}, // D02.2 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b01000011, 10'b1100010101, 2'b11}, // D03.2 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b01000011, 10'b1100010101, 2'b01}, // D03.2 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b01000100, 10'b1101010101, 2'b01}, // D04.2 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b01000100, 10'b0010100101, 2'b11}, // D04.2 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b01000101, 10'b1010010101, 2'b11}, // D05.2 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b01000101, 10'b1010010101, 2'b01}, // D05.2 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b01000110, 10'b0110010101, 2'b11}, // D06.2 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b01000110, 10'b0110010101, 2'b01}, // D06.2 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b01000111, 10'b1110000101, 2'b11}, // D07.2 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b01000111, 10'b0001110101, 2'b01}, // D07.2 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b01001000, 10'b1110010101, 2'b01}, // D08.2 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b01001000, 10'b0001100101, 2'b11}, // D08.2 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b01001001, 10'b1001010101, 2'b11}, // D09.2 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b01001001, 10'b1001010101, 2'b01}, // D09.2 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b01001010, 10'b0101010101, 2'b11}, // D10.2 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b01001010, 10'b0101010101, 2'b01}, // D10.2 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b01001011, 10'b1101000101, 2'b11}, // D11.2 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b01001011, 10'b1101000101, 2'b01}, // D11.2 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b01001100, 10'b0011010101, 2'b11}, // D12.2 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b01001100, 10'b0011010101, 2'b01}, // D12.2 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b01001101, 10'b1011000101, 2'b11}, // D13.2 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b01001101, 10'b1011000101, 2'b01}, // D13.2 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b01001110, 10'b0111000101, 2'b11}, // D14.2 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b01001110, 10'b0111000101, 2'b01}, // D14.2 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b01001111, 10'b0101110101, 2'b01}, // D15.2 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b01001111, 10'b1010000101, 2'b11}, // D15.2 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b01010000, 10'b0110110101, 2'b01}, // D16.2 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b01010000, 10'b1001000101, 2'b11}, // D16.2 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b01010001, 10'b1000110101, 2'b11}, // D17.2 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b01010001, 10'b1000110101, 2'b01}, // D17.2 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b01010010, 10'b0100110101, 2'b11}, // D18.2 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b01010010, 10'b0100110101, 2'b01}, // D18.2 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b01010011, 10'b1100100101, 2'b11}, // D19.2 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b01010011, 10'b1100100101, 2'b01}, // D19.2 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b01010100, 10'b0010110101, 2'b11}, // D20.2 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b01010100, 10'b0010110101, 2'b01}, // D20.2 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b01010101, 10'b1010100101, 2'b11}, // D21.2 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b01010101, 10'b1010100101, 2'b01}, // D21.2 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b01010110, 10'b0110100101, 2'b11}, // D22.2 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b01010110, 10'b0110100101, 2'b01}, // D22.2 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b01010111, 10'b1110100101, 2'b01}, // D23.2 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b01010111, 10'b0001010101, 2'b11}, // D23.2 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b01011000, 10'b1100110101, 2'b01}, // D24.2 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b01011000, 10'b0011000101, 2'b11}, // D24.2 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b01011001, 10'b1001100101, 2'b11}, // D25.2 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b01011001, 10'b1001100101, 2'b01}, // D25.2 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b01011010, 10'b0101100101, 2'b11}, // D26.2 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b01011010, 10'b0101100101, 2'b01}, // D26.2 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b01011011, 10'b1101100101, 2'b01}, // D27.2 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b01011011, 10'b0010010101, 2'b11}, // D27.2 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b01011100, 10'b0011100101, 2'b11}, // D28.2 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b01011100, 10'b0011100101, 2'b01}, // D28.2 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b01011101, 10'b1011100101, 2'b01}, // D29.2 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b01011101, 10'b0100010101, 2'b11}, // D29.2 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b01011110, 10'b0111100101, 2'b01}, // D30.2 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b01011110, 10'b1000010101, 2'b11}, // D30.2 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b01011111, 10'b1010110101, 2'b01}, // D31.2 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b01011111, 10'b0101000101, 2'b11}, // D31.2 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b01100000, 10'b1001110011, 2'b01}, // D00.3 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b01100000, 10'b0110001100, 2'b11}, // D00.3 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b01100001, 10'b0111010011, 2'b01}, // D01.3 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b01100001, 10'b1000101100, 2'b11}, // D01.3 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b01100010, 10'b1011010011, 2'b01}, // D02.3 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b01100010, 10'b0100101100, 2'b11}, // D02.3 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b01100011, 10'b1100011100, 2'b11}, // D03.3 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b01100011, 10'b1100010011, 2'b01}, // D03.3 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b01100100, 10'b1101010011, 2'b01}, // D04.3 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b01100100, 10'b0010101100, 2'b11}, // D04.3 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b01100101, 10'b1010011100, 2'b11}, // D05.3 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b01100101, 10'b1010010011, 2'b01}, // D05.3 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b01100110, 10'b0110011100, 2'b11}, // D06.3 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b01100110, 10'b0110010011, 2'b01}, // D06.3 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b01100111, 10'b1110001100, 2'b11}, // D07.3 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b01100111, 10'b0001110011, 2'b01}, // D07.3 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b01101000, 10'b1110010011, 2'b01}, // D08.3 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b01101000, 10'b0001101100, 2'b11}, // D08.3 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b01101001, 10'b1001011100, 2'b11}, // D09.3 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b01101001, 10'b1001010011, 2'b01}, // D09.3 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b01101010, 10'b0101011100, 2'b11}, // D10.3 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b01101010, 10'b0101010011, 2'b01}, // D10.3 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b01101011, 10'b1101001100, 2'b11}, // D11.3 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b01101011, 10'b1101000011, 2'b01}, // D11.3 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b01101100, 10'b0011011100, 2'b11}, // D12.3 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b01101100, 10'b0011010011, 2'b01}, // D12.3 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b01101101, 10'b1011001100, 2'b11}, // D13.3 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b01101101, 10'b1011000011, 2'b01}, // D13.3 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b01101110, 10'b0111001100, 2'b11}, // D14.3 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b01101110, 10'b0111000011, 2'b01}, // D14.3 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b01101111, 10'b0101110011, 2'b01}, // D15.3 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b01101111, 10'b1010001100, 2'b11}, // D15.3 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b01110000, 10'b0110110011, 2'b01}, // D16.3 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b01110000, 10'b1001001100, 2'b11}, // D16.3 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b01110001, 10'b1000111100, 2'b11}, // D17.3 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b01110001, 10'b1000110011, 2'b01}, // D17.3 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b01110010, 10'b0100111100, 2'b11}, // D18.3 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b01110010, 10'b0100110011, 2'b01}, // D18.3 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b01110011, 10'b1100101100, 2'b11}, // D19.3 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b01110011, 10'b1100100011, 2'b01}, // D19.3 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b01110100, 10'b0010111100, 2'b11}, // D20.3 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b01110100, 10'b0010110011, 2'b01}, // D20.3 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b01110101, 10'b1010101100, 2'b11}, // D21.3 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b01110101, 10'b1010100011, 2'b01}, // D21.3 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b01110110, 10'b0110101100, 2'b11}, // D22.3 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b01110110, 10'b0110100011, 2'b01}, // D22.3 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b01110111, 10'b1110100011, 2'b01}, // D23.3 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b01110111, 10'b0001011100, 2'b11}, // D23.3 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b01111000, 10'b1100110011, 2'b01}, // D24.3 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b01111000, 10'b0011001100, 2'b11}, // D24.3 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b01111001, 10'b1001101100, 2'b11}, // D25.3 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b01111001, 10'b1001100011, 2'b01}, // D25.3 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b01111010, 10'b0101101100, 2'b11}, // D26.3 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b01111010, 10'b0101100011, 2'b01}, // D26.3 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b01111011, 10'b1101100011, 2'b01}, // D27.3 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b01111011, 10'b0010011100, 2'b11}, // D27.3 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b01111100, 10'b0011101100, 2'b11}, // D28.3 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b01111100, 10'b0011100011, 2'b01}, // D28.3 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b01111101, 10'b1011100011, 2'b01}, // D29.3 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b01111101, 10'b0100011100, 2'b11}, // D29.3 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b01111110, 10'b0111100011, 2'b01}, // D30.3 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b01111110, 10'b1000011100, 2'b11}, // D30.3 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b01111111, 10'b1010110011, 2'b01}, // D31.3 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b01111111, 10'b0101001100, 2'b11}, // D31.3 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b10000000, 10'b1001110010, 2'b11}, // D00.4 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b10000000, 10'b0110001101, 2'b01}, // D00.4 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b10000001, 10'b0111010010, 2'b11}, // D01.4 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b10000001, 10'b1000101101, 2'b01}, // D01.4 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b10000010, 10'b1011010010, 2'b11}, // D02.4 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b10000010, 10'b0100101101, 2'b01}, // D02.4 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b10000011, 10'b1100011101, 2'b01}, // D03.4 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b10000011, 10'b1100010010, 2'b11}, // D03.4 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b10000100, 10'b1101010010, 2'b11}, // D04.4 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b10000100, 10'b0010101101, 2'b01}, // D04.4 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b10000101, 10'b1010011101, 2'b01}, // D05.4 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b10000101, 10'b1010010010, 2'b11}, // D05.4 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b10000110, 10'b0110011101, 2'b01}, // D06.4 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b10000110, 10'b0110010010, 2'b11}, // D06.4 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b10000111, 10'b1110001101, 2'b01}, // D07.4 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b10000111, 10'b0001110010, 2'b11}, // D07.4 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b10001000, 10'b1110010010, 2'b11}, // D08.4 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b10001000, 10'b0001101101, 2'b01}, // D08.4 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b10001001, 10'b1001011101, 2'b01}, // D09.4 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b10001001, 10'b1001010010, 2'b11}, // D09.4 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b10001010, 10'b0101011101, 2'b01}, // D10.4 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b10001010, 10'b0101010010, 2'b11}, // D10.4 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b10001011, 10'b1101001101, 2'b01}, // D11.4 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b10001011, 10'b1101000010, 2'b11}, // D11.4 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b10001100, 10'b0011011101, 2'b01}, // D12.4 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b10001100, 10'b0011010010, 2'b11}, // D12.4 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b10001101, 10'b1011001101, 2'b01}, // D13.4 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b10001101, 10'b1011000010, 2'b11}, // D13.4 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b10001110, 10'b0111001101, 2'b01}, // D14.4 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b10001110, 10'b0111000010, 2'b11}, // D14.4 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b10001111, 10'b0101110010, 2'b11}, // D15.4 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b10001111, 10'b1010001101, 2'b01}, // D15.4 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b10010000, 10'b0110110010, 2'b11}, // D16.4 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b10010000, 10'b1001001101, 2'b01}, // D16.4 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b10010001, 10'b1000111101, 2'b01}, // D17.4 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b10010001, 10'b1000110010, 2'b11}, // D17.4 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b10010010, 10'b0100111101, 2'b01}, // D18.4 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b10010010, 10'b0100110010, 2'b11}, // D18.4 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b10010011, 10'b1100101101, 2'b01}, // D19.4 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b10010011, 10'b1100100010, 2'b11}, // D19.4 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b10010100, 10'b0010111101, 2'b01}, // D20.4 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b10010100, 10'b0010110010, 2'b11}, // D20.4 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b10010101, 10'b1010101101, 2'b01}, // D21.4 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b10010101, 10'b1010100010, 2'b11}, // D21.4 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b10010110, 10'b0110101101, 2'b01}, // D22.4 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b10010110, 10'b0110100010, 2'b11}, // D22.4 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b10010111, 10'b1110100010, 2'b11}, // D23.4 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b10010111, 10'b0001011101, 2'b01}, // D23.4 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b10011000, 10'b1100110010, 2'b11}, // D24.4 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b10011000, 10'b0011001101, 2'b01}, // D24.4 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b10011001, 10'b1001101101, 2'b01}, // D25.4 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b10011001, 10'b1001100010, 2'b11}, // D25.4 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b10011010, 10'b0101101101, 2'b01}, // D26.4 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b10011010, 10'b0101100010, 2'b11}, // D26.4 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b10011011, 10'b1101100010, 2'b11}, // D27.4 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b10011011, 10'b0010011101, 2'b01}, // D27.4 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b10011100, 10'b0011101101, 2'b01}, // D28.4 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b10011100, 10'b0011100010, 2'b11}, // D28.4 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b10011101, 10'b1011100010, 2'b11}, // D29.4 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b10011101, 10'b0100011101, 2'b01}, // D29.4 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b10011110, 10'b0111100010, 2'b11}, // D30.4 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b10011110, 10'b1000011101, 2'b01}, // D30.4 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b10011111, 10'b1010110010, 2'b11}, // D31.4 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b10011111, 10'b0101001101, 2'b01}, // D31.4 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b10100000, 10'b1001111010, 2'b01}, // D00.5 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b10100000, 10'b0110001010, 2'b11}, // D00.5 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b10100001, 10'b0111011010, 2'b01}, // D01.5 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b10100001, 10'b1000101010, 2'b11}, // D01.5 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b10100010, 10'b1011011010, 2'b01}, // D02.5 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b10100010, 10'b0100101010, 2'b11}, // D02.5 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b10100011, 10'b1100011010, 2'b11}, // D03.5 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b10100011, 10'b1100011010, 2'b01}, // D03.5 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b10100100, 10'b1101011010, 2'b01}, // D04.5 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b10100100, 10'b0010101010, 2'b11}, // D04.5 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b10100101, 10'b1010011010, 2'b11}, // D05.5 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b10100101, 10'b1010011010, 2'b01}, // D05.5 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b10100110, 10'b0110011010, 2'b11}, // D06.5 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b10100110, 10'b0110011010, 2'b01}, // D06.5 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b10100111, 10'b1110001010, 2'b11}, // D07.5 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b10100111, 10'b0001111010, 2'b01}, // D07.5 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b10101000, 10'b1110011010, 2'b01}, // D08.5 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b10101000, 10'b0001101010, 2'b11}, // D08.5 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b10101001, 10'b1001011010, 2'b11}, // D09.5 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b10101001, 10'b1001011010, 2'b01}, // D09.5 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b10101010, 10'b0101011010, 2'b11}, // D10.5 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b10101010, 10'b0101011010, 2'b01}, // D10.5 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b10101011, 10'b1101001010, 2'b11}, // D11.5 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b10101011, 10'b1101001010, 2'b01}, // D11.5 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b10101100, 10'b0011011010, 2'b11}, // D12.5 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b10101100, 10'b0011011010, 2'b01}, // D12.5 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b10101101, 10'b1011001010, 2'b11}, // D13.5 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b10101101, 10'b1011001010, 2'b01}, // D13.5 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b10101110, 10'b0111001010, 2'b11}, // D14.5 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b10101110, 10'b0111001010, 2'b01}, // D14.5 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b10101111, 10'b0101111010, 2'b01}, // D15.5 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b10101111, 10'b1010001010, 2'b11}, // D15.5 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b10110000, 10'b0110111010, 2'b01}, // D16.5 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b10110000, 10'b1001001010, 2'b11}, // D16.5 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b10110001, 10'b1000111010, 2'b11}, // D17.5 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b10110001, 10'b1000111010, 2'b01}, // D17.5 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b10110010, 10'b0100111010, 2'b11}, // D18.5 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b10110010, 10'b0100111010, 2'b01}, // D18.5 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b10110011, 10'b1100101010, 2'b11}, // D19.5 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b10110011, 10'b1100101010, 2'b01}, // D19.5 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b10110100, 10'b0010111010, 2'b11}, // D20.5 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b10110100, 10'b0010111010, 2'b01}, // D20.5 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b10110101, 10'b1010101010, 2'b11}, // D21.5 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b10110101, 10'b1010101010, 2'b01}, // D21.5 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b10110110, 10'b0110101010, 2'b11}, // D22.5 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b10110110, 10'b0110101010, 2'b01}, // D22.5 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b10110111, 10'b1110101010, 2'b01}, // D23.5 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b10110111, 10'b0001011010, 2'b11}, // D23.5 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b10111000, 10'b1100111010, 2'b01}, // D24.5 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b10111000, 10'b0011001010, 2'b11}, // D24.5 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b10111001, 10'b1001101010, 2'b11}, // D25.5 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b10111001, 10'b1001101010, 2'b01}, // D25.5 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b10111010, 10'b0101101010, 2'b11}, // D26.5 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b10111010, 10'b0101101010, 2'b01}, // D26.5 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b10111011, 10'b1101101010, 2'b01}, // D27.5 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b10111011, 10'b0010011010, 2'b11}, // D27.5 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b10111100, 10'b0011101010, 2'b11}, // D28.5 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b10111100, 10'b0011101010, 2'b01}, // D28.5 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b10111101, 10'b1011101010, 2'b01}, // D29.5 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b10111101, 10'b0100011010, 2'b11}, // D29.5 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b10111110, 10'b0111101010, 2'b01}, // D30.5 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b10111110, 10'b1000011010, 2'b11}, // D30.5 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b10111111, 10'b1010111010, 2'b01}, // D31.5 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b10111111, 10'b0101001010, 2'b11}, // D31.5 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b11000000, 10'b1001110110, 2'b01}, // D00.6 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b11000000, 10'b0110000110, 2'b11}, // D00.6 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b11000001, 10'b0111010110, 2'b01}, // D01.6 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b11000001, 10'b1000100110, 2'b11}, // D01.6 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b11000010, 10'b1011010110, 2'b01}, // D02.6 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b11000010, 10'b0100100110, 2'b11}, // D02.6 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b11000011, 10'b1100010110, 2'b11}, // D03.6 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b11000011, 10'b1100010110, 2'b01}, // D03.6 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b11000100, 10'b1101010110, 2'b01}, // D04.6 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b11000100, 10'b0010100110, 2'b11}, // D04.6 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b11000101, 10'b1010010110, 2'b11}, // D05.6 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b11000101, 10'b1010010110, 2'b01}, // D05.6 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b11000110, 10'b0110010110, 2'b11}, // D06.6 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b11000110, 10'b0110010110, 2'b01}, // D06.6 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b11000111, 10'b1110000110, 2'b11}, // D07.6 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b11000111, 10'b0001110110, 2'b01}, // D07.6 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b11001000, 10'b1110010110, 2'b01}, // D08.6 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b11001000, 10'b0001100110, 2'b11}, // D08.6 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b11001001, 10'b1001010110, 2'b11}, // D09.6 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b11001001, 10'b1001010110, 2'b01}, // D09.6 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b11001010, 10'b0101010110, 2'b11}, // D10.6 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b11001010, 10'b0101010110, 2'b01}, // D10.6 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b11001011, 10'b1101000110, 2'b11}, // D11.6 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b11001011, 10'b1101000110, 2'b01}, // D11.6 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b11001100, 10'b0011010110, 2'b11}, // D12.6 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b11001100, 10'b0011010110, 2'b01}, // D12.6 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b11001101, 10'b1011000110, 2'b11}, // D13.6 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b11001101, 10'b1011000110, 2'b01}, // D13.6 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b11001110, 10'b0111000110, 2'b11}, // D14.6 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b11001110, 10'b0111000110, 2'b01}, // D14.6 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b11001111, 10'b0101110110, 2'b01}, // D15.6 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b11001111, 10'b1010000110, 2'b11}, // D15.6 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b11010000, 10'b0110110110, 2'b01}, // D16.6 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b11010000, 10'b1001000110, 2'b11}, // D16.6 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b11010001, 10'b1000110110, 2'b11}, // D17.6 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b11010001, 10'b1000110110, 2'b01}, // D17.6 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b11010010, 10'b0100110110, 2'b11}, // D18.6 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b11010010, 10'b0100110110, 2'b01}, // D18.6 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b11010011, 10'b1100100110, 2'b11}, // D19.6 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b11010011, 10'b1100100110, 2'b01}, // D19.6 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b11010100, 10'b0010110110, 2'b11}, // D20.6 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b11010100, 10'b0010110110, 2'b01}, // D20.6 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b11010101, 10'b1010100110, 2'b11}, // D21.6 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b11010101, 10'b1010100110, 2'b01}, // D21.6 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b11010110, 10'b0110100110, 2'b11}, // D22.6 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b11010110, 10'b0110100110, 2'b01}, // D22.6 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b11010111, 10'b1110100110, 2'b01}, // D23.6 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b11010111, 10'b0001010110, 2'b11}, // D23.6 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b11011000, 10'b1100110110, 2'b01}, // D24.6 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b11011000, 10'b0011000110, 2'b11}, // D24.6 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b11011001, 10'b1001100110, 2'b11}, // D25.6 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b11011001, 10'b1001100110, 2'b01}, // D25.6 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b11011010, 10'b0101100110, 2'b11}, // D26.6 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b11011010, 10'b0101100110, 2'b01}, // D26.6 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b11011011, 10'b1101100110, 2'b01}, // D27.6 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b11011011, 10'b0010010110, 2'b11}, // D27.6 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b11011100, 10'b0011100110, 2'b11}, // D28.6 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b11011100, 10'b0011100110, 2'b01}, // D28.6 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b11011101, 10'b1011100110, 2'b01}, // D29.6 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b11011101, 10'b0100010110, 2'b11}, // D29.6 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b11011110, 10'b0111100110, 2'b01}, // D30.6 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b11011110, 10'b1000010110, 2'b11}, // D30.6 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b11011111, 10'b1010110110, 2'b01}, // D31.6 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b11011111, 10'b0101000110, 2'b11}, // D31.6 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b11100000, 10'b1001110001, 2'b11}, // D00.7 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b11100000, 10'b0110001110, 2'b01}, // D00.7 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b11100001, 10'b0111010001, 2'b11}, // D01.7 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b11100001, 10'b1000101110, 2'b01}, // D01.7 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b11100010, 10'b1011010001, 2'b11}, // D02.7 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b11100010, 10'b0100101110, 2'b01}, // D02.7 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b11100011, 10'b1100011110, 2'b01}, // D03.7 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b11100011, 10'b1100010001, 2'b11}, // D03.7 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b11100100, 10'b1101010001, 2'b11}, // D04.7 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b11100100, 10'b0010101110, 2'b01}, // D04.7 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b11100101, 10'b1010011110, 2'b01}, // D05.7 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b11100101, 10'b1010010001, 2'b11}, // D05.7 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b11100110, 10'b0110011110, 2'b01}, // D06.7 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b11100110, 10'b0110010001, 2'b11}, // D06.7 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b11100111, 10'b1110001110, 2'b01}, // D07.7 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b11100111, 10'b0001110001, 2'b11}, // D07.7 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b11101000, 10'b1110010001, 2'b11}, // D08.7 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b11101000, 10'b0001101110, 2'b01}, // D08.7 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b11101001, 10'b1001011110, 2'b01}, // D09.7 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b11101001, 10'b1001010001, 2'b11}, // D09.7 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b11101010, 10'b0101011110, 2'b01}, // D10.7 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b11101010, 10'b0101010001, 2'b11}, // D10.7 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b11101011, 10'b1101001110, 2'b01}, // D11.7 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b11101011, 10'b1101001000, 2'b11}, // D11.7 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b11101100, 10'b0011011110, 2'b01}, // D12.7 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b11101100, 10'b0011010001, 2'b11}, // D12.7 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b11101101, 10'b1011001110, 2'b01}, // D13.7 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b11101101, 10'b1011001000, 2'b11}, // D13.7 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b11101110, 10'b0111001110, 2'b01}, // D14.7 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b11101110, 10'b0111001000, 2'b11}, // D14.7 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b11101111, 10'b0101110001, 2'b11}, // D15.7 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b11101111, 10'b1010001110, 2'b01}, // D15.7 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b11110000, 10'b0110110001, 2'b11}, // D16.7 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b11110000, 10'b1001001110, 2'b01}, // D16.7 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b11110001, 10'b1000110111, 2'b01}, // D17.7 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b11110001, 10'b1000110001, 2'b11}, // D17.7 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b11110010, 10'b0100110111, 2'b01}, // D18.7 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b11110010, 10'b0100110001, 2'b11}, // D18.7 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b11110011, 10'b1100101110, 2'b01}, // D19.7 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b11110011, 10'b1100100001, 2'b11}, // D19.7 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b11110100, 10'b0010110111, 2'b01}, // D20.7 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b11110100, 10'b0010110001, 2'b11}, // D20.7 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b11110101, 10'b1010101110, 2'b01}, // D21.7 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b11110101, 10'b1010100001, 2'b11}, // D21.7 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b11110110, 10'b0110101110, 2'b01}, // D22.7 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b11110110, 10'b0110100001, 2'b11}, // D22.7 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b11110111, 10'b1110100001, 2'b11}, // D23.7 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b11110111, 10'b0001011110, 2'b01}, // D23.7 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b11111000, 10'b1100110001, 2'b11}, // D24.7 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b11111000, 10'b0011001110, 2'b01}, // D24.7 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b11111001, 10'b1001101110, 2'b01}, // D25.7 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b11111001, 10'b1001100001, 2'b11}, // D25.7 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b11111010, 10'b0101101110, 2'b01}, // D26.7 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b11111010, 10'b0101100001, 2'b11}, // D26.7 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b11111011, 10'b1101100001, 2'b11}, // D27.7 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b11111011, 10'b0010011110, 2'b01}, // D27.7 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b11111100, 10'b0011101110, 2'b01}, // D28.7 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b11111100, 10'b0011100001, 2'b11}, // D28.7 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b11111101, 10'b1011100001, 2'b11}, // D29.7 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b11111101, 10'b0100011110, 2'b01}, // D29.7 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b11111110, 10'b0111100001, 2'b11}, // D30.7 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b11111110, 10'b1000011110, 2'b01}, // D30.7 (RD = +1)
   {1'b0, 1'b0, 2'b11, 8'b11111111, 10'b1010110001, 2'b11}, // D31.7 (RD = -1)
   {1'b0, 1'b0, 2'b01, 8'b11111111, 10'b0101001110, 2'b01}, // D31.7 (RD = +1)
   {1'b1, 1'b1, 2'b11, 8'b00000000, 10'b1001110100, 2'b11}, // ?
   {1'b1, 1'b1, 2'b01, 8'b00000000, 10'b0110001011, 2'b01}, // ?
   {1'b1, 1'b1, 2'b11, 8'b00000001, 10'b0111010100, 2'b11}, // ?
   {1'b1, 1'b1, 2'b01, 8'b00000001, 10'b1000101011, 2'b01}, // ?
   {1'b1, 1'b1, 2'b11, 8'b00000010, 10'b1011010100, 2'b11}, // ?
   {1'b1, 1'b1, 2'b01, 8'b00000010, 10'b0100101011, 2'b01}, // ?
   {1'b1, 1'b1, 2'b11, 8'b00000011, 10'b1100011011, 2'b01}, // ?
   {1'b1, 1'b1, 2'b01, 8'b00000011, 10'b1100010100, 2'b11}, // ?
   {1'b1, 1'b1, 2'b11, 8'b00000100, 10'b1101010100, 2'b11}, // ?
   {1'b1, 1'b1, 2'b01, 8'b00000100, 10'b0010101011, 2'b01}, // ?
   {1'b1, 1'b1, 2'b11, 8'b00000101, 10'b1010011011, 2'b01}, // ?
   {1'b1, 1'b1, 2'b01, 8'b00000101, 10'b1010010100, 2'b11}, // ?
   {1'b1, 1'b1, 2'b11, 8'b00000110, 10'b0110011011, 2'b01}, // ?
   {1'b1, 1'b1, 2'b01, 8'b00000110, 10'b0110010100, 2'b11}, // ?
   {1'b1, 1'b1, 2'b11, 8'b00000111, 10'b1110001011, 2'b01}, // ?
   {1'b1, 1'b1, 2'b01, 8'b00000111, 10'b0001110100, 2'b11}, // ?
   {1'b1, 1'b1, 2'b11, 8'b00001000, 10'b1110010100, 2'b11}, // ?
   {1'b1, 1'b1, 2'b01, 8'b00001000, 10'b0001101011, 2'b01}, // ?
   {1'b1, 1'b1, 2'b11, 8'b00001001, 10'b1001011011, 2'b01}, // ?
   {1'b1, 1'b1, 2'b01, 8'b00001001, 10'b1001010100, 2'b11}, // ?
   {1'b1, 1'b1, 2'b11, 8'b00001010, 10'b0101011011, 2'b01}, // ?
   {1'b1, 1'b1, 2'b01, 8'b00001010, 10'b0101010100, 2'b11}, // ?
   {1'b1, 1'b1, 2'b11, 8'b00001011, 10'b1101001011, 2'b01}, // ?
   {1'b1, 1'b1, 2'b01, 8'b00001011, 10'b1101000100, 2'b11}, // ?
   {1'b1, 1'b1, 2'b11, 8'b00001100, 10'b0011011011, 2'b01}, // ?
   {1'b1, 1'b1, 2'b01, 8'b00001100, 10'b0011010100, 2'b11}, // ?
   {1'b1, 1'b1, 2'b11, 8'b00001101, 10'b1011001011, 2'b01}, // ?
   {1'b1, 1'b1, 2'b01, 8'b00001101, 10'b1011000100, 2'b11}, // ?
   {1'b1, 1'b1, 2'b11, 8'b00001110, 10'b0111001011, 2'b01}, // ?
   {1'b1, 1'b1, 2'b01, 8'b00001110, 10'b0111000100, 2'b11}, // ?
   {1'b1, 1'b1, 2'b11, 8'b00001111, 10'b0101110100, 2'b11}, // ?
   {1'b1, 1'b1, 2'b01, 8'b00001111, 10'b1010001011, 2'b01}, // ?
   {1'b1, 1'b1, 2'b11, 8'b00010000, 10'b0110110100, 2'b11}, // ?
   {1'b1, 1'b1, 2'b01, 8'b00010000, 10'b1001001011, 2'b01}, // ?
   {1'b1, 1'b1, 2'b11, 8'b00010001, 10'b1000111011, 2'b01}, // ?
   {1'b1, 1'b1, 2'b01, 8'b00010001, 10'b1000110100, 2'b11}, // ?
   {1'b1, 1'b1, 2'b11, 8'b00010010, 10'b0100111011, 2'b01}, // ?
   {1'b1, 1'b1, 2'b01, 8'b00010010, 10'b0100110100, 2'b11}, // ?
   {1'b1, 1'b1, 2'b11, 8'b00010011, 10'b1100101011, 2'b01}, // ?
   {1'b1, 1'b1, 2'b01, 8'b00010011, 10'b1100100100, 2'b11}, // ?
   {1'b1, 1'b1, 2'b11, 8'b00010100, 10'b0010111011, 2'b01}, // ?
   {1'b1, 1'b1, 2'b01, 8'b00010100, 10'b0010110100, 2'b11}, // ?
   {1'b1, 1'b1, 2'b11, 8'b00010101, 10'b1010101011, 2'b01}, // ?
   {1'b1, 1'b1, 2'b01, 8'b00010101, 10'b1010100100, 2'b11}, // ?
   {1'b1, 1'b1, 2'b11, 8'b00010110, 10'b0110101011, 2'b01}, // ?
   {1'b1, 1'b1, 2'b01, 8'b00010110, 10'b0110100100, 2'b11}, // ?
   {1'b1, 1'b1, 2'b11, 8'b00010111, 10'b1110100100, 2'b11}, // ?
   {1'b1, 1'b1, 2'b01, 8'b00010111, 10'b0001011011, 2'b01}, // ?
   {1'b1, 1'b1, 2'b11, 8'b00011000, 10'b1100110100, 2'b11}, // ?
   {1'b1, 1'b1, 2'b01, 8'b00011000, 10'b0011001011, 2'b01}, // ?
   {1'b1, 1'b1, 2'b11, 8'b00011001, 10'b1001101011, 2'b01}, // ?
   {1'b1, 1'b1, 2'b01, 8'b00011001, 10'b1001100100, 2'b11}, // ?
   {1'b1, 1'b1, 2'b11, 8'b00011010, 10'b0101101011, 2'b01}, // ?
   {1'b1, 1'b1, 2'b01, 8'b00011010, 10'b0101100100, 2'b11}, // ?
   {1'b1, 1'b1, 2'b11, 8'b00011011, 10'b1101100100, 2'b11}, // ?
   {1'b1, 1'b1, 2'b01, 8'b00011011, 10'b0010011011, 2'b01}, // ?
   {1'b0, 1'b1, 2'b11, 8'b00011100, 10'b0011110100, 2'b11}, // K28.0 (RD = -1)
   {1'b0, 1'b1, 2'b01, 8'b00011100, 10'b1100001011, 2'b01}, // K28.0 (RD = +1)
   {1'b1, 1'b1, 2'b11, 8'b00011101, 10'b1011100100, 2'b11}, // ?
   {1'b1, 1'b1, 2'b01, 8'b00011101, 10'b0100011011, 2'b01}, // ?
   {1'b1, 1'b1, 2'b11, 8'b00011110, 10'b0111100100, 2'b11}, // ?
   {1'b1, 1'b1, 2'b01, 8'b00011110, 10'b1000011011, 2'b01}, // ?
   {1'b1, 1'b1, 2'b11, 8'b00011111, 10'b1010110100, 2'b11}, // ?
   {1'b1, 1'b1, 2'b01, 8'b00011111, 10'b0101001011, 2'b01}, // ?
   {1'b1, 1'b1, 2'b11, 8'b00100000, 10'b1001111001, 2'b01}, // ?
   {1'b1, 1'b1, 2'b01, 8'b00100000, 10'b0110001001, 2'b11}, // ?
   {1'b1, 1'b1, 2'b11, 8'b00100001, 10'b0111011001, 2'b01}, // ?
   {1'b1, 1'b1, 2'b01, 8'b00100001, 10'b1000101001, 2'b11}, // ?
   {1'b1, 1'b1, 2'b11, 8'b00100010, 10'b1011011001, 2'b01}, // ?
   {1'b1, 1'b1, 2'b01, 8'b00100010, 10'b0100101001, 2'b11}, // ?
   {1'b1, 1'b1, 2'b11, 8'b00100011, 10'b1100011001, 2'b11}, // ?
   {1'b1, 1'b1, 2'b01, 8'b00100011, 10'b1100011001, 2'b01}, // ?
   {1'b1, 1'b1, 2'b11, 8'b00100100, 10'b1101011001, 2'b01}, // ?
   {1'b1, 1'b1, 2'b01, 8'b00100100, 10'b0010101001, 2'b11}, // ?
   {1'b1, 1'b1, 2'b11, 8'b00100101, 10'b1010011001, 2'b11}, // ?
   {1'b1, 1'b1, 2'b01, 8'b00100101, 10'b1010011001, 2'b01}, // ?
   {1'b1, 1'b1, 2'b11, 8'b00100110, 10'b0110011001, 2'b11}, // ?
   {1'b1, 1'b1, 2'b01, 8'b00100110, 10'b0110011001, 2'b01}, // ?
   {1'b1, 1'b1, 2'b11, 8'b00100111, 10'b1110001001, 2'b11}, // ?
   {1'b1, 1'b1, 2'b01, 8'b00100111, 10'b0001111001, 2'b01}, // ?
   {1'b1, 1'b1, 2'b11, 8'b00101000, 10'b1110011001, 2'b01}, // ?
   {1'b1, 1'b1, 2'b01, 8'b00101000, 10'b0001101001, 2'b11}, // ?
   {1'b1, 1'b1, 2'b11, 8'b00101001, 10'b1001011001, 2'b11}, // ?
   {1'b1, 1'b1, 2'b01, 8'b00101001, 10'b1001011001, 2'b01}, // ?
   {1'b1, 1'b1, 2'b11, 8'b00101010, 10'b0101011001, 2'b11}, // ?
   {1'b1, 1'b1, 2'b01, 8'b00101010, 10'b0101011001, 2'b01}, // ?
   {1'b1, 1'b1, 2'b11, 8'b00101011, 10'b1101001001, 2'b11}, // ?
   {1'b1, 1'b1, 2'b01, 8'b00101011, 10'b1101001001, 2'b01}, // ?
   {1'b1, 1'b1, 2'b11, 8'b00101100, 10'b0011011001, 2'b11}, // ?
   {1'b1, 1'b1, 2'b01, 8'b00101100, 10'b0011011001, 2'b01}, // ?
   {1'b1, 1'b1, 2'b11, 8'b00101101, 10'b1011001001, 2'b11}, // ?
   {1'b1, 1'b1, 2'b01, 8'b00101101, 10'b1011001001, 2'b01}, // ?
   {1'b1, 1'b1, 2'b11, 8'b00101110, 10'b0111001001, 2'b11}, // ?
   {1'b1, 1'b1, 2'b01, 8'b00101110, 10'b0111001001, 2'b01}, // ?
   {1'b1, 1'b1, 2'b11, 8'b00101111, 10'b0101111001, 2'b01}, // ?
   {1'b1, 1'b1, 2'b01, 8'b00101111, 10'b1010001001, 2'b11}, // ?
   {1'b1, 1'b1, 2'b11, 8'b00110000, 10'b0110111001, 2'b01}, // ?
   {1'b1, 1'b1, 2'b01, 8'b00110000, 10'b1001001001, 2'b11}, // ?
   {1'b1, 1'b1, 2'b11, 8'b00110001, 10'b1000111001, 2'b11}, // ?
   {1'b1, 1'b1, 2'b01, 8'b00110001, 10'b1000111001, 2'b01}, // ?
   {1'b1, 1'b1, 2'b11, 8'b00110010, 10'b0100111001, 2'b11}, // ?
   {1'b1, 1'b1, 2'b01, 8'b00110010, 10'b0100111001, 2'b01}, // ?
   {1'b1, 1'b1, 2'b11, 8'b00110011, 10'b1100101001, 2'b11}, // ?
   {1'b1, 1'b1, 2'b01, 8'b00110011, 10'b1100101001, 2'b01}, // ?
   {1'b1, 1'b1, 2'b11, 8'b00110100, 10'b0010111001, 2'b11}, // ?
   {1'b1, 1'b1, 2'b01, 8'b00110100, 10'b0010111001, 2'b01}, // ?
   {1'b1, 1'b1, 2'b11, 8'b00110101, 10'b1010101001, 2'b11}, // ?
   {1'b1, 1'b1, 2'b01, 8'b00110101, 10'b1010101001, 2'b01}, // ?
   {1'b1, 1'b1, 2'b11, 8'b00110110, 10'b0110101001, 2'b11}, // ?
   {1'b1, 1'b1, 2'b01, 8'b00110110, 10'b0110101001, 2'b01}, // ?
   {1'b1, 1'b1, 2'b11, 8'b00110111, 10'b1110101001, 2'b01}, // ?
   {1'b1, 1'b1, 2'b01, 8'b00110111, 10'b0001011001, 2'b11}, // ?
   {1'b1, 1'b1, 2'b11, 8'b00111000, 10'b1100111001, 2'b01}, // ?
   {1'b1, 1'b1, 2'b01, 8'b00111000, 10'b0011001001, 2'b11}, // ?
   {1'b1, 1'b1, 2'b11, 8'b00111001, 10'b1001101001, 2'b11}, // ?
   {1'b1, 1'b1, 2'b01, 8'b00111001, 10'b1001101001, 2'b01}, // ?
   {1'b1, 1'b1, 2'b11, 8'b00111010, 10'b0101101001, 2'b11}, // ?
   {1'b1, 1'b1, 2'b01, 8'b00111010, 10'b0101101001, 2'b01}, // ?
   {1'b1, 1'b1, 2'b11, 8'b00111011, 10'b1101101001, 2'b01}, // ?
   {1'b1, 1'b1, 2'b01, 8'b00111011, 10'b0010011001, 2'b11}, // ?
   {1'b0, 1'b1, 2'b11, 8'b00111100, 10'b0011111001, 2'b01}, // K28.1 (RD = -1)
   {1'b0, 1'b1, 2'b01, 8'b00111100, 10'b1100000110, 2'b11}, // K28.1 (RD = +1)
   {1'b1, 1'b1, 2'b11, 8'b00111101, 10'b1011101001, 2'b01}, // ?
   {1'b1, 1'b1, 2'b01, 8'b00111101, 10'b0100011001, 2'b11}, // ?
   {1'b1, 1'b1, 2'b11, 8'b00111110, 10'b0111101001, 2'b01}, // ?
   {1'b1, 1'b1, 2'b01, 8'b00111110, 10'b1000011001, 2'b11}, // ?
   {1'b1, 1'b1, 2'b11, 8'b00111111, 10'b1010111001, 2'b01}, // ?
   {1'b1, 1'b1, 2'b01, 8'b00111111, 10'b0101001001, 2'b11}, // ?
   {1'b1, 1'b1, 2'b11, 8'b01000000, 10'b1001110101, 2'b01}, // ?
   {1'b1, 1'b1, 2'b01, 8'b01000000, 10'b0110000101, 2'b11}, // ?
   {1'b1, 1'b1, 2'b11, 8'b01000001, 10'b0111010101, 2'b01}, // ?
   {1'b1, 1'b1, 2'b01, 8'b01000001, 10'b1000100101, 2'b11}, // ?
   {1'b1, 1'b1, 2'b11, 8'b01000010, 10'b1011010101, 2'b01}, // ?
   {1'b1, 1'b1, 2'b01, 8'b01000010, 10'b0100100101, 2'b11}, // ?
   {1'b1, 1'b1, 2'b11, 8'b01000011, 10'b1100010101, 2'b11}, // ?
   {1'b1, 1'b1, 2'b01, 8'b01000011, 10'b1100010101, 2'b01}, // ?
   {1'b1, 1'b1, 2'b11, 8'b01000100, 10'b1101010101, 2'b01}, // ?
   {1'b1, 1'b1, 2'b01, 8'b01000100, 10'b0010100101, 2'b11}, // ?
   {1'b1, 1'b1, 2'b11, 8'b01000101, 10'b1010010101, 2'b11}, // ?
   {1'b1, 1'b1, 2'b01, 8'b01000101, 10'b1010010101, 2'b01}, // ?
   {1'b1, 1'b1, 2'b11, 8'b01000110, 10'b0110010101, 2'b11}, // ?
   {1'b1, 1'b1, 2'b01, 8'b01000110, 10'b0110010101, 2'b01}, // ?
   {1'b1, 1'b1, 2'b11, 8'b01000111, 10'b1110000101, 2'b11}, // ?
   {1'b1, 1'b1, 2'b01, 8'b01000111, 10'b0001110101, 2'b01}, // ?
   {1'b1, 1'b1, 2'b11, 8'b01001000, 10'b1110010101, 2'b01}, // ?
   {1'b1, 1'b1, 2'b01, 8'b01001000, 10'b0001100101, 2'b11}, // ?
   {1'b1, 1'b1, 2'b11, 8'b01001001, 10'b1001010101, 2'b11}, // ?
   {1'b1, 1'b1, 2'b01, 8'b01001001, 10'b1001010101, 2'b01}, // ?
   {1'b1, 1'b1, 2'b11, 8'b01001010, 10'b0101010101, 2'b11}, // ?
   {1'b1, 1'b1, 2'b01, 8'b01001010, 10'b0101010101, 2'b01}, // ?
   {1'b1, 1'b1, 2'b11, 8'b01001011, 10'b1101000101, 2'b11}, // ?
   {1'b1, 1'b1, 2'b01, 8'b01001011, 10'b1101000101, 2'b01}, // ?
   {1'b1, 1'b1, 2'b11, 8'b01001100, 10'b0011010101, 2'b11}, // ?
   {1'b1, 1'b1, 2'b01, 8'b01001100, 10'b0011010101, 2'b01}, // ?
   {1'b1, 1'b1, 2'b11, 8'b01001101, 10'b1011000101, 2'b11}, // ?
   {1'b1, 1'b1, 2'b01, 8'b01001101, 10'b1011000101, 2'b01}, // ?
   {1'b1, 1'b1, 2'b11, 8'b01001110, 10'b0111000101, 2'b11}, // ?
   {1'b1, 1'b1, 2'b01, 8'b01001110, 10'b0111000101, 2'b01}, // ?
   {1'b1, 1'b1, 2'b11, 8'b01001111, 10'b0101110101, 2'b01}, // ?
   {1'b1, 1'b1, 2'b01, 8'b01001111, 10'b1010000101, 2'b11}, // ?
   {1'b1, 1'b1, 2'b11, 8'b01010000, 10'b0110110101, 2'b01}, // ?
   {1'b1, 1'b1, 2'b01, 8'b01010000, 10'b1001000101, 2'b11}, // ?
   {1'b1, 1'b1, 2'b11, 8'b01010001, 10'b1000110101, 2'b11}, // ?
   {1'b1, 1'b1, 2'b01, 8'b01010001, 10'b1000110101, 2'b01}, // ?
   {1'b1, 1'b1, 2'b11, 8'b01010010, 10'b0100110101, 2'b11}, // ?
   {1'b1, 1'b1, 2'b01, 8'b01010010, 10'b0100110101, 2'b01}, // ?
   {1'b1, 1'b1, 2'b11, 8'b01010011, 10'b1100100101, 2'b11}, // ?
   {1'b1, 1'b1, 2'b01, 8'b01010011, 10'b1100100101, 2'b01}, // ?
   {1'b1, 1'b1, 2'b11, 8'b01010100, 10'b0010110101, 2'b11}, // ?
   {1'b1, 1'b1, 2'b01, 8'b01010100, 10'b0010110101, 2'b01}, // ?
   {1'b1, 1'b1, 2'b11, 8'b01010101, 10'b1010100101, 2'b11}, // ?
   {1'b1, 1'b1, 2'b01, 8'b01010101, 10'b1010100101, 2'b01}, // ?
   {1'b1, 1'b1, 2'b11, 8'b01010110, 10'b0110100101, 2'b11}, // ?
   {1'b1, 1'b1, 2'b01, 8'b01010110, 10'b0110100101, 2'b01}, // ?
   {1'b1, 1'b1, 2'b11, 8'b01010111, 10'b1110100101, 2'b01}, // ?
   {1'b1, 1'b1, 2'b01, 8'b01010111, 10'b0001010101, 2'b11}, // ?
   {1'b1, 1'b1, 2'b11, 8'b01011000, 10'b1100110101, 2'b01}, // ?
   {1'b1, 1'b1, 2'b01, 8'b01011000, 10'b0011000101, 2'b11}, // ?
   {1'b1, 1'b1, 2'b11, 8'b01011001, 10'b1001100101, 2'b11}, // ?
   {1'b1, 1'b1, 2'b01, 8'b01011001, 10'b1001100101, 2'b01}, // ?
   {1'b1, 1'b1, 2'b11, 8'b01011010, 10'b0101100101, 2'b11}, // ?
   {1'b1, 1'b1, 2'b01, 8'b01011010, 10'b0101100101, 2'b01}, // ?
   {1'b1, 1'b1, 2'b11, 8'b01011011, 10'b1101100101, 2'b01}, // ?
   {1'b1, 1'b1, 2'b01, 8'b01011011, 10'b0010010101, 2'b11}, // ?
   {1'b0, 1'b1, 2'b11, 8'b01011100, 10'b0011110101, 2'b01}, // K28.2 (RD = -1)
   {1'b0, 1'b1, 2'b01, 8'b01011100, 10'b1100001010, 2'b11}, // K28.2 (RD = +1)
   {1'b1, 1'b1, 2'b11, 8'b01011101, 10'b1011100101, 2'b01}, // ?
   {1'b1, 1'b1, 2'b01, 8'b01011101, 10'b0100010101, 2'b11}, // ?
   {1'b1, 1'b1, 2'b11, 8'b01011110, 10'b0111100101, 2'b01}, // ?
   {1'b1, 1'b1, 2'b01, 8'b01011110, 10'b1000010101, 2'b11}, // ?
   {1'b1, 1'b1, 2'b11, 8'b01011111, 10'b1010110101, 2'b01}, // ?
   {1'b1, 1'b1, 2'b01, 8'b01011111, 10'b0101000101, 2'b11}, // ?
   {1'b1, 1'b1, 2'b11, 8'b01100000, 10'b1001110011, 2'b01}, // ?
   {1'b1, 1'b1, 2'b01, 8'b01100000, 10'b0110001100, 2'b11}, // ?
   {1'b1, 1'b1, 2'b11, 8'b01100001, 10'b0111010011, 2'b01}, // ?
   {1'b1, 1'b1, 2'b01, 8'b01100001, 10'b1000101100, 2'b11}, // ?
   {1'b1, 1'b1, 2'b11, 8'b01100010, 10'b1011010011, 2'b01}, // ?
   {1'b1, 1'b1, 2'b01, 8'b01100010, 10'b0100101100, 2'b11}, // ?
   {1'b1, 1'b1, 2'b11, 8'b01100011, 10'b1100011100, 2'b11}, // ?
   {1'b1, 1'b1, 2'b01, 8'b01100011, 10'b1100010011, 2'b01}, // ?
   {1'b1, 1'b1, 2'b11, 8'b01100100, 10'b1101010011, 2'b01}, // ?
   {1'b1, 1'b1, 2'b01, 8'b01100100, 10'b0010101100, 2'b11}, // ?
   {1'b1, 1'b1, 2'b11, 8'b01100101, 10'b1010011100, 2'b11}, // ?
   {1'b1, 1'b1, 2'b01, 8'b01100101, 10'b1010010011, 2'b01}, // ?
   {1'b1, 1'b1, 2'b11, 8'b01100110, 10'b0110011100, 2'b11}, // ?
   {1'b1, 1'b1, 2'b01, 8'b01100110, 10'b0110010011, 2'b01}, // ?
   {1'b1, 1'b1, 2'b11, 8'b01100111, 10'b1110001100, 2'b11}, // ?
   {1'b1, 1'b1, 2'b01, 8'b01100111, 10'b0001110011, 2'b01}, // ?
   {1'b1, 1'b1, 2'b11, 8'b01101000, 10'b1110010011, 2'b01}, // ?
   {1'b1, 1'b1, 2'b01, 8'b01101000, 10'b0001101100, 2'b11}, // ?
   {1'b1, 1'b1, 2'b11, 8'b01101001, 10'b1001011100, 2'b11}, // ?
   {1'b1, 1'b1, 2'b01, 8'b01101001, 10'b1001010011, 2'b01}, // ?
   {1'b1, 1'b1, 2'b11, 8'b01101010, 10'b0101011100, 2'b11}, // ?
   {1'b1, 1'b1, 2'b01, 8'b01101010, 10'b0101010011, 2'b01}, // ?
   {1'b1, 1'b1, 2'b11, 8'b01101011, 10'b1101001100, 2'b11}, // ?
   {1'b1, 1'b1, 2'b01, 8'b01101011, 10'b1101000011, 2'b01}, // ?
   {1'b1, 1'b1, 2'b11, 8'b01101100, 10'b0011011100, 2'b11}, // ?
   {1'b1, 1'b1, 2'b01, 8'b01101100, 10'b0011010011, 2'b01}, // ?
   {1'b1, 1'b1, 2'b11, 8'b01101101, 10'b1011001100, 2'b11}, // ?
   {1'b1, 1'b1, 2'b01, 8'b01101101, 10'b1011000011, 2'b01}, // ?
   {1'b1, 1'b1, 2'b11, 8'b01101110, 10'b0111001100, 2'b11}, // ?
   {1'b1, 1'b1, 2'b01, 8'b01101110, 10'b0111000011, 2'b01}, // ?
   {1'b1, 1'b1, 2'b11, 8'b01101111, 10'b0101110011, 2'b01}, // ?
   {1'b1, 1'b1, 2'b01, 8'b01101111, 10'b1010001100, 2'b11}, // ?
   {1'b1, 1'b1, 2'b11, 8'b01110000, 10'b0110110011, 2'b01}, // ?
   {1'b1, 1'b1, 2'b01, 8'b01110000, 10'b1001001100, 2'b11}, // ?
   {1'b1, 1'b1, 2'b11, 8'b01110001, 10'b1000111100, 2'b11}, // ?
   {1'b1, 1'b1, 2'b01, 8'b01110001, 10'b1000110011, 2'b01}, // ?
   {1'b1, 1'b1, 2'b11, 8'b01110010, 10'b0100111100, 2'b11}, // ?
   {1'b1, 1'b1, 2'b01, 8'b01110010, 10'b0100110011, 2'b01}, // ?
   {1'b1, 1'b1, 2'b11, 8'b01110011, 10'b1100101100, 2'b11}, // ?
   {1'b1, 1'b1, 2'b01, 8'b01110011, 10'b1100100011, 2'b01}, // ?
   {1'b1, 1'b1, 2'b11, 8'b01110100, 10'b0010111100, 2'b11}, // ?
   {1'b1, 1'b1, 2'b01, 8'b01110100, 10'b0010110011, 2'b01}, // ?
   {1'b1, 1'b1, 2'b11, 8'b01110101, 10'b1010101100, 2'b11}, // ?
   {1'b1, 1'b1, 2'b01, 8'b01110101, 10'b1010100011, 2'b01}, // ?
   {1'b1, 1'b1, 2'b11, 8'b01110110, 10'b0110101100, 2'b11}, // ?
   {1'b1, 1'b1, 2'b01, 8'b01110110, 10'b0110100011, 2'b01}, // ?
   {1'b1, 1'b1, 2'b11, 8'b01110111, 10'b1110100011, 2'b01}, // ?
   {1'b1, 1'b1, 2'b01, 8'b01110111, 10'b0001011100, 2'b11}, // ?
   {1'b1, 1'b1, 2'b11, 8'b01111000, 10'b1100110011, 2'b01}, // ?
   {1'b1, 1'b1, 2'b01, 8'b01111000, 10'b0011001100, 2'b11}, // ?
   {1'b1, 1'b1, 2'b11, 8'b01111001, 10'b1001101100, 2'b11}, // ?
   {1'b1, 1'b1, 2'b01, 8'b01111001, 10'b1001100011, 2'b01}, // ?
   {1'b1, 1'b1, 2'b11, 8'b01111010, 10'b0101101100, 2'b11}, // ?
   {1'b1, 1'b1, 2'b01, 8'b01111010, 10'b0101100011, 2'b01}, // ?
   {1'b1, 1'b1, 2'b11, 8'b01111011, 10'b1101100011, 2'b01}, // ?
   {1'b1, 1'b1, 2'b01, 8'b01111011, 10'b0010011100, 2'b11}, // ?
   {1'b0, 1'b1, 2'b11, 8'b01111100, 10'b0011110011, 2'b01}, // K28.3 (RD = -1)
   {1'b0, 1'b1, 2'b01, 8'b01111100, 10'b1100001100, 2'b11}, // K28.3 (RD = +1)
   {1'b1, 1'b1, 2'b11, 8'b01111101, 10'b1011100011, 2'b01}, // ?
   {1'b1, 1'b1, 2'b01, 8'b01111101, 10'b0100011100, 2'b11}, // ?
   {1'b1, 1'b1, 2'b11, 8'b01111110, 10'b0111100011, 2'b01}, // ?
   {1'b1, 1'b1, 2'b01, 8'b01111110, 10'b1000011100, 2'b11}, // ?
   {1'b1, 1'b1, 2'b11, 8'b01111111, 10'b1010110011, 2'b01}, // ?
   {1'b1, 1'b1, 2'b01, 8'b01111111, 10'b0101001100, 2'b11}, // ?
   {1'b1, 1'b1, 2'b11, 8'b10000000, 10'b1001110010, 2'b11}, // ?
   {1'b1, 1'b1, 2'b01, 8'b10000000, 10'b0110001101, 2'b01}, // ?
   {1'b1, 1'b1, 2'b11, 8'b10000001, 10'b0111010010, 2'b11}, // ?
   {1'b1, 1'b1, 2'b01, 8'b10000001, 10'b1000101101, 2'b01}, // ?
   {1'b1, 1'b1, 2'b11, 8'b10000010, 10'b1011010010, 2'b11}, // ?
   {1'b1, 1'b1, 2'b01, 8'b10000010, 10'b0100101101, 2'b01}, // ?
   {1'b1, 1'b1, 2'b11, 8'b10000011, 10'b1100011101, 2'b01}, // ?
   {1'b1, 1'b1, 2'b01, 8'b10000011, 10'b1100010010, 2'b11}, // ?
   {1'b1, 1'b1, 2'b11, 8'b10000100, 10'b1101010010, 2'b11}, // ?
   {1'b1, 1'b1, 2'b01, 8'b10000100, 10'b0010101101, 2'b01}, // ?
   {1'b1, 1'b1, 2'b11, 8'b10000101, 10'b1010011101, 2'b01}, // ?
   {1'b1, 1'b1, 2'b01, 8'b10000101, 10'b1010010010, 2'b11}, // ?
   {1'b1, 1'b1, 2'b11, 8'b10000110, 10'b0110011101, 2'b01}, // ?
   {1'b1, 1'b1, 2'b01, 8'b10000110, 10'b0110010010, 2'b11}, // ?
   {1'b1, 1'b1, 2'b11, 8'b10000111, 10'b1110001101, 2'b01}, // ?
   {1'b1, 1'b1, 2'b01, 8'b10000111, 10'b0001110010, 2'b11}, // ?
   {1'b1, 1'b1, 2'b11, 8'b10001000, 10'b1110010010, 2'b11}, // ?
   {1'b1, 1'b1, 2'b01, 8'b10001000, 10'b0001101101, 2'b01}, // ?
   {1'b1, 1'b1, 2'b11, 8'b10001001, 10'b1001011101, 2'b01}, // ?
   {1'b1, 1'b1, 2'b01, 8'b10001001, 10'b1001010010, 2'b11}, // ?
   {1'b1, 1'b1, 2'b11, 8'b10001010, 10'b0101011101, 2'b01}, // ?
   {1'b1, 1'b1, 2'b01, 8'b10001010, 10'b0101010010, 2'b11}, // ?
   {1'b1, 1'b1, 2'b11, 8'b10001011, 10'b1101001101, 2'b01}, // ?
   {1'b1, 1'b1, 2'b01, 8'b10001011, 10'b1101000010, 2'b11}, // ?
   {1'b1, 1'b1, 2'b11, 8'b10001100, 10'b0011011101, 2'b01}, // ?
   {1'b1, 1'b1, 2'b01, 8'b10001100, 10'b0011010010, 2'b11}, // ?
   {1'b1, 1'b1, 2'b11, 8'b10001101, 10'b1011001101, 2'b01}, // ?
   {1'b1, 1'b1, 2'b01, 8'b10001101, 10'b1011000010, 2'b11}, // ?
   {1'b1, 1'b1, 2'b11, 8'b10001110, 10'b0111001101, 2'b01}, // ?
   {1'b1, 1'b1, 2'b01, 8'b10001110, 10'b0111000010, 2'b11}, // ?
   {1'b1, 1'b1, 2'b11, 8'b10001111, 10'b0101110010, 2'b11}, // ?
   {1'b1, 1'b1, 2'b01, 8'b10001111, 10'b1010001101, 2'b01}, // ?
   {1'b1, 1'b1, 2'b11, 8'b10010000, 10'b0110110010, 2'b11}, // ?
   {1'b1, 1'b1, 2'b01, 8'b10010000, 10'b1001001101, 2'b01}, // ?
   {1'b1, 1'b1, 2'b11, 8'b10010001, 10'b1000111101, 2'b01}, // ?
   {1'b1, 1'b1, 2'b01, 8'b10010001, 10'b1000110010, 2'b11}, // ?
   {1'b1, 1'b1, 2'b11, 8'b10010010, 10'b0100111101, 2'b01}, // ?
   {1'b1, 1'b1, 2'b01, 8'b10010010, 10'b0100110010, 2'b11}, // ?
   {1'b1, 1'b1, 2'b11, 8'b10010011, 10'b1100101101, 2'b01}, // ?
   {1'b1, 1'b1, 2'b01, 8'b10010011, 10'b1100100010, 2'b11}, // ?
   {1'b1, 1'b1, 2'b11, 8'b10010100, 10'b0010111101, 2'b01}, // ?
   {1'b1, 1'b1, 2'b01, 8'b10010100, 10'b0010110010, 2'b11}, // ?
   {1'b1, 1'b1, 2'b11, 8'b10010101, 10'b1010101101, 2'b01}, // ?
   {1'b1, 1'b1, 2'b01, 8'b10010101, 10'b1010100010, 2'b11}, // ?
   {1'b1, 1'b1, 2'b11, 8'b10010110, 10'b0110101101, 2'b01}, // ?
   {1'b1, 1'b1, 2'b01, 8'b10010110, 10'b0110100010, 2'b11}, // ?
   {1'b1, 1'b1, 2'b11, 8'b10010111, 10'b1110100010, 2'b11}, // ?
   {1'b1, 1'b1, 2'b01, 8'b10010111, 10'b0001011101, 2'b01}, // ?
   {1'b1, 1'b1, 2'b11, 8'b10011000, 10'b1100110010, 2'b11}, // ?
   {1'b1, 1'b1, 2'b01, 8'b10011000, 10'b0011001101, 2'b01}, // ?
   {1'b1, 1'b1, 2'b11, 8'b10011001, 10'b1001101101, 2'b01}, // ?
   {1'b1, 1'b1, 2'b01, 8'b10011001, 10'b1001100010, 2'b11}, // ?
   {1'b1, 1'b1, 2'b11, 8'b10011010, 10'b0101101101, 2'b01}, // ?
   {1'b1, 1'b1, 2'b01, 8'b10011010, 10'b0101100010, 2'b11}, // ?
   {1'b1, 1'b1, 2'b11, 8'b10011011, 10'b1101100010, 2'b11}, // ?
   {1'b1, 1'b1, 2'b01, 8'b10011011, 10'b0010011101, 2'b01}, // ?
   {1'b0, 1'b1, 2'b11, 8'b10011100, 10'b0011110010, 2'b11}, // K28.4 (RD = -1)
   {1'b0, 1'b1, 2'b01, 8'b10011100, 10'b1100001101, 2'b01}, // K28.4 (RD = +1)
   {1'b1, 1'b1, 2'b11, 8'b10011101, 10'b1011100010, 2'b11}, // ?
   {1'b1, 1'b1, 2'b01, 8'b10011101, 10'b0100011101, 2'b01}, // ?
   {1'b1, 1'b1, 2'b11, 8'b10011110, 10'b0111100010, 2'b11}, // ?
   {1'b1, 1'b1, 2'b01, 8'b10011110, 10'b1000011101, 2'b01}, // ?
   {1'b1, 1'b1, 2'b11, 8'b10011111, 10'b1010110010, 2'b11}, // ?
   {1'b1, 1'b1, 2'b01, 8'b10011111, 10'b0101001101, 2'b01}, // ?
   {1'b1, 1'b1, 2'b11, 8'b10100000, 10'b1001111010, 2'b01}, // ?
   {1'b1, 1'b1, 2'b01, 8'b10100000, 10'b0110001010, 2'b11}, // ?
   {1'b1, 1'b1, 2'b11, 8'b10100001, 10'b0111011010, 2'b01}, // ?
   {1'b1, 1'b1, 2'b01, 8'b10100001, 10'b1000101010, 2'b11}, // ?
   {1'b1, 1'b1, 2'b11, 8'b10100010, 10'b1011011010, 2'b01}, // ?
   {1'b1, 1'b1, 2'b01, 8'b10100010, 10'b0100101010, 2'b11}, // ?
   {1'b1, 1'b1, 2'b11, 8'b10100011, 10'b1100011010, 2'b11}, // ?
   {1'b1, 1'b1, 2'b01, 8'b10100011, 10'b1100011010, 2'b01}, // ?
   {1'b1, 1'b1, 2'b11, 8'b10100100, 10'b1101011010, 2'b01}, // ?
   {1'b1, 1'b1, 2'b01, 8'b10100100, 10'b0010101010, 2'b11}, // ?
   {1'b1, 1'b1, 2'b11, 8'b10100101, 10'b1010011010, 2'b11}, // ?
   {1'b1, 1'b1, 2'b01, 8'b10100101, 10'b1010011010, 2'b01}, // ?
   {1'b1, 1'b1, 2'b11, 8'b10100110, 10'b0110011010, 2'b11}, // ?
   {1'b1, 1'b1, 2'b01, 8'b10100110, 10'b0110011010, 2'b01}, // ?
   {1'b1, 1'b1, 2'b11, 8'b10100111, 10'b1110001010, 2'b11}, // ?
   {1'b1, 1'b1, 2'b01, 8'b10100111, 10'b0001111010, 2'b01}, // ?
   {1'b1, 1'b1, 2'b11, 8'b10101000, 10'b1110011010, 2'b01}, // ?
   {1'b1, 1'b1, 2'b01, 8'b10101000, 10'b0001101010, 2'b11}, // ?
   {1'b1, 1'b1, 2'b11, 8'b10101001, 10'b1001011010, 2'b11}, // ?
   {1'b1, 1'b1, 2'b01, 8'b10101001, 10'b1001011010, 2'b01}, // ?
   {1'b1, 1'b1, 2'b11, 8'b10101010, 10'b0101011010, 2'b11}, // ?
   {1'b1, 1'b1, 2'b01, 8'b10101010, 10'b0101011010, 2'b01}, // ?
   {1'b1, 1'b1, 2'b11, 8'b10101011, 10'b1101001010, 2'b11}, // ?
   {1'b1, 1'b1, 2'b01, 8'b10101011, 10'b1101001010, 2'b01}, // ?
   {1'b1, 1'b1, 2'b11, 8'b10101100, 10'b0011011010, 2'b11}, // ?
   {1'b1, 1'b1, 2'b01, 8'b10101100, 10'b0011011010, 2'b01}, // ?
   {1'b1, 1'b1, 2'b11, 8'b10101101, 10'b1011001010, 2'b11}, // ?
   {1'b1, 1'b1, 2'b01, 8'b10101101, 10'b1011001010, 2'b01}, // ?
   {1'b1, 1'b1, 2'b11, 8'b10101110, 10'b0111001010, 2'b11}, // ?
   {1'b1, 1'b1, 2'b01, 8'b10101110, 10'b0111001010, 2'b01}, // ?
   {1'b1, 1'b1, 2'b11, 8'b10101111, 10'b0101111010, 2'b01}, // ?
   {1'b1, 1'b1, 2'b01, 8'b10101111, 10'b1010001010, 2'b11}, // ?
   {1'b1, 1'b1, 2'b11, 8'b10110000, 10'b0110111010, 2'b01}, // ?
   {1'b1, 1'b1, 2'b01, 8'b10110000, 10'b1001001010, 2'b11}, // ?
   {1'b1, 1'b1, 2'b11, 8'b10110001, 10'b1000111010, 2'b11}, // ?
   {1'b1, 1'b1, 2'b01, 8'b10110001, 10'b1000111010, 2'b01}, // ?
   {1'b1, 1'b1, 2'b11, 8'b10110010, 10'b0100111010, 2'b11}, // ?
   {1'b1, 1'b1, 2'b01, 8'b10110010, 10'b0100111010, 2'b01}, // ?
   {1'b1, 1'b1, 2'b11, 8'b10110011, 10'b1100101010, 2'b11}, // ?
   {1'b1, 1'b1, 2'b01, 8'b10110011, 10'b1100101010, 2'b01}, // ?
   {1'b1, 1'b1, 2'b11, 8'b10110100, 10'b0010111010, 2'b11}, // ?
   {1'b1, 1'b1, 2'b01, 8'b10110100, 10'b0010111010, 2'b01}, // ?
   {1'b1, 1'b1, 2'b11, 8'b10110101, 10'b1010101010, 2'b11}, // ?
   {1'b1, 1'b1, 2'b01, 8'b10110101, 10'b1010101010, 2'b01}, // ?
   {1'b1, 1'b1, 2'b11, 8'b10110110, 10'b0110101010, 2'b11}, // ?
   {1'b1, 1'b1, 2'b01, 8'b10110110, 10'b0110101010, 2'b01}, // ?
   {1'b1, 1'b1, 2'b11, 8'b10110111, 10'b1110101010, 2'b01}, // ?
   {1'b1, 1'b1, 2'b01, 8'b10110111, 10'b0001011010, 2'b11}, // ?
   {1'b1, 1'b1, 2'b11, 8'b10111000, 10'b1100111010, 2'b01}, // ?
   {1'b1, 1'b1, 2'b01, 8'b10111000, 10'b0011001010, 2'b11}, // ?
   {1'b1, 1'b1, 2'b11, 8'b10111001, 10'b1001101010, 2'b11}, // ?
   {1'b1, 1'b1, 2'b01, 8'b10111001, 10'b1001101010, 2'b01}, // ?
   {1'b1, 1'b1, 2'b11, 8'b10111010, 10'b0101101010, 2'b11}, // ?
   {1'b1, 1'b1, 2'b01, 8'b10111010, 10'b0101101010, 2'b01}, // ?
   {1'b1, 1'b1, 2'b11, 8'b10111011, 10'b1101101010, 2'b01}, // ?
   {1'b1, 1'b1, 2'b01, 8'b10111011, 10'b0010011010, 2'b11}, // ?
   {1'b0, 1'b1, 2'b11, 8'b10111100, 10'b0011111010, 2'b01}, // K28.5 (RD = -1)
   {1'b0, 1'b1, 2'b01, 8'b10111100, 10'b1100000101, 2'b11}, // K28.5 (RD = +1)
   {1'b1, 1'b1, 2'b11, 8'b10111101, 10'b1011101010, 2'b01}, // ?
   {1'b1, 1'b1, 2'b01, 8'b10111101, 10'b0100011010, 2'b11}, // ?
   {1'b1, 1'b1, 2'b11, 8'b10111110, 10'b0111101010, 2'b01}, // ?
   {1'b1, 1'b1, 2'b01, 8'b10111110, 10'b1000011010, 2'b11}, // ?
   {1'b1, 1'b1, 2'b11, 8'b10111111, 10'b1010111010, 2'b01}, // ?
   {1'b1, 1'b1, 2'b01, 8'b10111111, 10'b0101001010, 2'b11}, // ?
   {1'b1, 1'b1, 2'b11, 8'b11000000, 10'b1001110110, 2'b01}, // ?
   {1'b1, 1'b1, 2'b01, 8'b11000000, 10'b0110000110, 2'b11}, // ?
   {1'b1, 1'b1, 2'b11, 8'b11000001, 10'b0111010110, 2'b01}, // ?
   {1'b1, 1'b1, 2'b01, 8'b11000001, 10'b1000100110, 2'b11}, // ?
   {1'b1, 1'b1, 2'b11, 8'b11000010, 10'b1011010110, 2'b01}, // ?
   {1'b1, 1'b1, 2'b01, 8'b11000010, 10'b0100100110, 2'b11}, // ?
   {1'b1, 1'b1, 2'b11, 8'b11000011, 10'b1100010110, 2'b11}, // ?
   {1'b1, 1'b1, 2'b01, 8'b11000011, 10'b1100010110, 2'b01}, // ?
   {1'b1, 1'b1, 2'b11, 8'b11000100, 10'b1101010110, 2'b01}, // ?
   {1'b1, 1'b1, 2'b01, 8'b11000100, 10'b0010100110, 2'b11}, // ?
   {1'b1, 1'b1, 2'b11, 8'b11000101, 10'b1010010110, 2'b11}, // ?
   {1'b1, 1'b1, 2'b01, 8'b11000101, 10'b1010010110, 2'b01}, // ?
   {1'b1, 1'b1, 2'b11, 8'b11000110, 10'b0110010110, 2'b11}, // ?
   {1'b1, 1'b1, 2'b01, 8'b11000110, 10'b0110010110, 2'b01}, // ?
   {1'b1, 1'b1, 2'b11, 8'b11000111, 10'b1110000110, 2'b11}, // ?
   {1'b1, 1'b1, 2'b01, 8'b11000111, 10'b0001110110, 2'b01}, // ?
   {1'b1, 1'b1, 2'b11, 8'b11001000, 10'b1110010110, 2'b01}, // ?
   {1'b1, 1'b1, 2'b01, 8'b11001000, 10'b0001100110, 2'b11}, // ?
   {1'b1, 1'b1, 2'b11, 8'b11001001, 10'b1001010110, 2'b11}, // ?
   {1'b1, 1'b1, 2'b01, 8'b11001001, 10'b1001010110, 2'b01}, // ?
   {1'b1, 1'b1, 2'b11, 8'b11001010, 10'b0101010110, 2'b11}, // ?
   {1'b1, 1'b1, 2'b01, 8'b11001010, 10'b0101010110, 2'b01}, // ?
   {1'b1, 1'b1, 2'b11, 8'b11001011, 10'b1101000110, 2'b11}, // ?
   {1'b1, 1'b1, 2'b01, 8'b11001011, 10'b1101000110, 2'b01}, // ?
   {1'b1, 1'b1, 2'b11, 8'b11001100, 10'b0011010110, 2'b11}, // ?
   {1'b1, 1'b1, 2'b01, 8'b11001100, 10'b0011010110, 2'b01}, // ?
   {1'b1, 1'b1, 2'b11, 8'b11001101, 10'b1011000110, 2'b11}, // ?
   {1'b1, 1'b1, 2'b01, 8'b11001101, 10'b1011000110, 2'b01}, // ?
   {1'b1, 1'b1, 2'b11, 8'b11001110, 10'b0111000110, 2'b11}, // ?
   {1'b1, 1'b1, 2'b01, 8'b11001110, 10'b0111000110, 2'b01}, // ?
   {1'b1, 1'b1, 2'b11, 8'b11001111, 10'b0101110110, 2'b01}, // ?
   {1'b1, 1'b1, 2'b01, 8'b11001111, 10'b1010000110, 2'b11}, // ?
   {1'b1, 1'b1, 2'b11, 8'b11010000, 10'b0110110110, 2'b01}, // ?
   {1'b1, 1'b1, 2'b01, 8'b11010000, 10'b1001000110, 2'b11}, // ?
   {1'b1, 1'b1, 2'b11, 8'b11010001, 10'b1000110110, 2'b11}, // ?
   {1'b1, 1'b1, 2'b01, 8'b11010001, 10'b1000110110, 2'b01}, // ?
   {1'b1, 1'b1, 2'b11, 8'b11010010, 10'b0100110110, 2'b11}, // ?
   {1'b1, 1'b1, 2'b01, 8'b11010010, 10'b0100110110, 2'b01}, // ?
   {1'b1, 1'b1, 2'b11, 8'b11010011, 10'b1100100110, 2'b11}, // ?
   {1'b1, 1'b1, 2'b01, 8'b11010011, 10'b1100100110, 2'b01}, // ?
   {1'b1, 1'b1, 2'b11, 8'b11010100, 10'b0010110110, 2'b11}, // ?
   {1'b1, 1'b1, 2'b01, 8'b11010100, 10'b0010110110, 2'b01}, // ?
   {1'b1, 1'b1, 2'b11, 8'b11010101, 10'b1010100110, 2'b11}, // ?
   {1'b1, 1'b1, 2'b01, 8'b11010101, 10'b1010100110, 2'b01}, // ?
   {1'b1, 1'b1, 2'b11, 8'b11010110, 10'b0110100110, 2'b11}, // ?
   {1'b1, 1'b1, 2'b01, 8'b11010110, 10'b0110100110, 2'b01}, // ?
   {1'b1, 1'b1, 2'b11, 8'b11010111, 10'b1110100110, 2'b01}, // ?
   {1'b1, 1'b1, 2'b01, 8'b11010111, 10'b0001010110, 2'b11}, // ?
   {1'b1, 1'b1, 2'b11, 8'b11011000, 10'b1100110110, 2'b01}, // ?
   {1'b1, 1'b1, 2'b01, 8'b11011000, 10'b0011000110, 2'b11}, // ?
   {1'b1, 1'b1, 2'b11, 8'b11011001, 10'b1001100110, 2'b11}, // ?
   {1'b1, 1'b1, 2'b01, 8'b11011001, 10'b1001100110, 2'b01}, // ?
   {1'b1, 1'b1, 2'b11, 8'b11011010, 10'b0101100110, 2'b11}, // ?
   {1'b1, 1'b1, 2'b01, 8'b11011010, 10'b0101100110, 2'b01}, // ?
   {1'b1, 1'b1, 2'b11, 8'b11011011, 10'b1101100110, 2'b01}, // ?
   {1'b1, 1'b1, 2'b01, 8'b11011011, 10'b0010010110, 2'b11}, // ?
   {1'b0, 1'b1, 2'b11, 8'b11011100, 10'b0011110110, 2'b01}, // K28.6 (RD = -1)
   {1'b0, 1'b1, 2'b01, 8'b11011100, 10'b1100001001, 2'b11}, // K28.6 (RD = +1)
   {1'b1, 1'b1, 2'b11, 8'b11011101, 10'b1011100110, 2'b01}, // ?
   {1'b1, 1'b1, 2'b01, 8'b11011101, 10'b0100010110, 2'b11}, // ?
   {1'b1, 1'b1, 2'b11, 8'b11011110, 10'b0111100110, 2'b01}, // ?
   {1'b1, 1'b1, 2'b01, 8'b11011110, 10'b1000010110, 2'b11}, // ?
   {1'b1, 1'b1, 2'b11, 8'b11011111, 10'b1010110110, 2'b01}, // ?
   {1'b1, 1'b1, 2'b01, 8'b11011111, 10'b0101000110, 2'b11}, // ?
   {1'b1, 1'b1, 2'b11, 8'b11100000, 10'b1001110001, 2'b11}, // ?
   {1'b1, 1'b1, 2'b01, 8'b11100000, 10'b0110001110, 2'b01}, // ?
   {1'b1, 1'b1, 2'b11, 8'b11100001, 10'b0111010001, 2'b11}, // ?
   {1'b1, 1'b1, 2'b01, 8'b11100001, 10'b1000101110, 2'b01}, // ?
   {1'b1, 1'b1, 2'b11, 8'b11100010, 10'b1011010001, 2'b11}, // ?
   {1'b1, 1'b1, 2'b01, 8'b11100010, 10'b0100101110, 2'b01}, // ?
   {1'b1, 1'b1, 2'b11, 8'b11100011, 10'b1100011110, 2'b01}, // ?
   {1'b1, 1'b1, 2'b01, 8'b11100011, 10'b1100010001, 2'b11}, // ?
   {1'b1, 1'b1, 2'b11, 8'b11100100, 10'b1101010001, 2'b11}, // ?
   {1'b1, 1'b1, 2'b01, 8'b11100100, 10'b0010101110, 2'b01}, // ?
   {1'b1, 1'b1, 2'b11, 8'b11100101, 10'b1010011110, 2'b01}, // ?
   {1'b1, 1'b1, 2'b01, 8'b11100101, 10'b1010010001, 2'b11}, // ?
   {1'b1, 1'b1, 2'b11, 8'b11100110, 10'b0110011110, 2'b01}, // ?
   {1'b1, 1'b1, 2'b01, 8'b11100110, 10'b0110010001, 2'b11}, // ?
   {1'b1, 1'b1, 2'b11, 8'b11100111, 10'b1110001110, 2'b01}, // ?
   {1'b1, 1'b1, 2'b01, 8'b11100111, 10'b0001110001, 2'b11}, // ?
   {1'b1, 1'b1, 2'b11, 8'b11101000, 10'b1110010001, 2'b11}, // ?
   {1'b1, 1'b1, 2'b01, 8'b11101000, 10'b0001101110, 2'b01}, // ?
   {1'b1, 1'b1, 2'b11, 8'b11101001, 10'b1001011110, 2'b01}, // ?
   {1'b1, 1'b1, 2'b01, 8'b11101001, 10'b1001010001, 2'b11}, // ?
   {1'b1, 1'b1, 2'b11, 8'b11101010, 10'b0101011110, 2'b01}, // ?
   {1'b1, 1'b1, 2'b01, 8'b11101010, 10'b0101010001, 2'b11}, // ?
   {1'b1, 1'b1, 2'b11, 8'b11101011, 10'b1101001110, 2'b01}, // ?
   {1'b1, 1'b1, 2'b01, 8'b11101011, 10'b1101001000, 2'b11}, // ?
   {1'b1, 1'b1, 2'b11, 8'b11101100, 10'b0011011110, 2'b01}, // ?
   {1'b1, 1'b1, 2'b01, 8'b11101100, 10'b0011010001, 2'b11}, // ?
   {1'b1, 1'b1, 2'b11, 8'b11101101, 10'b1011001110, 2'b01}, // ?
   {1'b1, 1'b1, 2'b01, 8'b11101101, 10'b1011001000, 2'b11}, // ?
   {1'b1, 1'b1, 2'b11, 8'b11101110, 10'b0111001110, 2'b01}, // ?
   {1'b1, 1'b1, 2'b01, 8'b11101110, 10'b0111001000, 2'b11}, // ?
   {1'b1, 1'b1, 2'b11, 8'b11101111, 10'b0101110001, 2'b11}, // ?
   {1'b1, 1'b1, 2'b01, 8'b11101111, 10'b1010001110, 2'b01}, // ?
   {1'b1, 1'b1, 2'b11, 8'b11110000, 10'b0110110001, 2'b11}, // ?
   {1'b1, 1'b1, 2'b01, 8'b11110000, 10'b1001001110, 2'b01}, // ?
   {1'b1, 1'b1, 2'b11, 8'b11110001, 10'b1000110111, 2'b01}, // ?
   {1'b1, 1'b1, 2'b01, 8'b11110001, 10'b1000110001, 2'b11}, // ?
   {1'b1, 1'b1, 2'b11, 8'b11110010, 10'b0100110111, 2'b01}, // ?
   {1'b1, 1'b1, 2'b01, 8'b11110010, 10'b0100110001, 2'b11}, // ?
   {1'b1, 1'b1, 2'b11, 8'b11110011, 10'b1100101110, 2'b01}, // ?
   {1'b1, 1'b1, 2'b01, 8'b11110011, 10'b1100100001, 2'b11}, // ?
   {1'b1, 1'b1, 2'b11, 8'b11110100, 10'b0010110111, 2'b01}, // ?
   {1'b1, 1'b1, 2'b01, 8'b11110100, 10'b0010110001, 2'b11}, // ?
   {1'b1, 1'b1, 2'b11, 8'b11110101, 10'b1010101110, 2'b01}, // ?
   {1'b1, 1'b1, 2'b01, 8'b11110101, 10'b1010100001, 2'b11}, // ?
   {1'b1, 1'b1, 2'b11, 8'b11110110, 10'b0110101110, 2'b01}, // ?
   {1'b1, 1'b1, 2'b01, 8'b11110110, 10'b0110100001, 2'b11}, // ?
   {1'b0, 1'b1, 2'b11, 8'b11110111, 10'b1110101000, 2'b11}, // K23.7 (RD = -1)
   {1'b0, 1'b1, 2'b01, 8'b11110111, 10'b0001010111, 2'b01}, // K23.7 (RD = +1)
   {1'b1, 1'b1, 2'b11, 8'b11111000, 10'b1100110001, 2'b11}, // ?
   {1'b1, 1'b1, 2'b01, 8'b11111000, 10'b0011001110, 2'b01}, // ?
   {1'b1, 1'b1, 2'b11, 8'b11111001, 10'b1001101110, 2'b01}, // ?
   {1'b1, 1'b1, 2'b01, 8'b11111001, 10'b1001100001, 2'b11}, // ?
   {1'b1, 1'b1, 2'b11, 8'b11111010, 10'b0101101110, 2'b01}, // ?
   {1'b1, 1'b1, 2'b01, 8'b11111010, 10'b0101100001, 2'b11}, // ?
   {1'b0, 1'b1, 2'b11, 8'b11111011, 10'b1101101000, 2'b11}, // K27.7 (RD = -1)
   {1'b0, 1'b1, 2'b01, 8'b11111011, 10'b0010010111, 2'b01}, // K27.7 (RD = +1)
   {1'b0, 1'b1, 2'b11, 8'b11111100, 10'b0011111000, 2'b11}, // K28.7 (RD = -1)
   {1'b0, 1'b1, 2'b01, 8'b11111100, 10'b1100000111, 2'b01}, // K28.7 (RD = +1)
   {1'b0, 1'b1, 2'b11, 8'b11111101, 10'b1011101000, 2'b11}, // K29.7 (RD = -1)
   {1'b0, 1'b1, 2'b01, 8'b11111101, 10'b0100010111, 2'b01}, // K29.7 (RD = +1)
   {1'b0, 1'b1, 2'b11, 8'b11111110, 10'b0111101000, 2'b11}, // K30.7 (RD = -1)
   {1'b0, 1'b1, 2'b01, 8'b11111110, 10'b1000010111, 2'b01}, // K30.7 (RD = +1)
   {1'b1, 1'b1, 2'b11, 8'b11111111, 10'b1010110001, 2'b11}, // ?
   {1'b1, 1'b1, 2'b01, 8'b11111111, 10'b0101001110, 2'b01}  // ?
  };

  string enc_byte_name [1024] = '{
    "D00.0 (RD = -1)",
    "D00.0 (RD = +1)",
    "D01.0 (RD = -1)",
    "D01.0 (RD = +1)",
    "D02.0 (RD = -1)",
    "D02.0 (RD = +1)",
    "D03.0 (RD = -1)",
    "D03.0 (RD = +1)",
    "D04.0 (RD = -1)",
    "D04.0 (RD = +1)",
    "D05.0 (RD = -1)",
    "D05.0 (RD = +1)",
    "D06.0 (RD = -1)",
    "D06.0 (RD = +1)",
    "D07.0 (RD = -1)",
    "D07.0 (RD = +1)",
    "D08.0 (RD = -1)",
    "D08.0 (RD = +1)",
    "D09.0 (RD = -1)",
    "D09.0 (RD = +1)",
    "D10.0 (RD = -1)",
    "D10.0 (RD = +1)",
    "D11.0 (RD = -1)",
    "D11.0 (RD = +1)",
    "D12.0 (RD = -1)",
    "D12.0 (RD = +1)",
    "D13.0 (RD = -1)",
    "D13.0 (RD = +1)",
    "D14.0 (RD = -1)",
    "D14.0 (RD = +1)",
    "D15.0 (RD = -1)",
    "D15.0 (RD = +1)",
    "D16.0 (RD = -1)",
    "D16.0 (RD = +1)",
    "D17.0 (RD = -1)",
    "D17.0 (RD = +1)",
    "D18.0 (RD = -1)",
    "D18.0 (RD = +1)",
    "D19.0 (RD = -1)",
    "D19.0 (RD = +1)",
    "D20.0 (RD = -1)",
    "D20.0 (RD = +1)",
    "D21.0 (RD = -1)",
    "D21.0 (RD = +1)",
    "D22.0 (RD = -1)",
    "D22.0 (RD = +1)",
    "D23.0 (RD = -1)",
    "D23.0 (RD = +1)",
    "D24.0 (RD = -1)",
    "D24.0 (RD = +1)",
    "D25.0 (RD = -1)",
    "D25.0 (RD = +1)",
    "D26.0 (RD = -1)",
    "D26.0 (RD = +1)",
    "D27.0 (RD = -1)",
    "D27.0 (RD = +1)",
    "D28.0 (RD = -1)",
    "D28.0 (RD = +1)",
    "D29.0 (RD = -1)",
    "D29.0 (RD = +1)",
    "D30.0 (RD = -1)",
    "D30.0 (RD = +1)",
    "D31.0 (RD = -1)",
    "D31.0 (RD = +1)",
    "D00.1 (RD = -1)",
    "D00.1 (RD = +1)",
    "D01.1 (RD = -1)",
    "D01.1 (RD = +1)",
    "D02.1 (RD = -1)",
    "D02.1 (RD = +1)",
    "D03.1 (RD = -1)",
    "D03.1 (RD = +1)",
    "D04.1 (RD = -1)",
    "D04.1 (RD = +1)",
    "D05.1 (RD = -1)",
    "D05.1 (RD = +1)",
    "D06.1 (RD = -1)",
    "D06.1 (RD = +1)",
    "D07.1 (RD = -1)",
    "D07.1 (RD = +1)",
    "D08.1 (RD = -1)",
    "D08.1 (RD = +1)",
    "D09.1 (RD = -1)",
    "D09.1 (RD = +1)",
    "D10.1 (RD = -1)",
    "D10.1 (RD = +1)",
    "D11.1 (RD = -1)",
    "D11.1 (RD = +1)",
    "D12.1 (RD = -1)",
    "D12.1 (RD = +1)",
    "D13.1 (RD = -1)",
    "D13.1 (RD = +1)",
    "D14.1 (RD = -1)",
    "D14.1 (RD = +1)",
    "D15.1 (RD = -1)",
    "D15.1 (RD = +1)",
    "D16.1 (RD = -1)",
    "D16.1 (RD = +1)",
    "D17.1 (RD = -1)",
    "D17.1 (RD = +1)",
    "D18.1 (RD = -1)",
    "D18.1 (RD = +1)",
    "D19.1 (RD = -1)",
    "D19.1 (RD = +1)",
    "D20.1 (RD = -1)",
    "D20.1 (RD = +1)",
    "D21.1 (RD = -1)",
    "D21.1 (RD = +1)",
    "D22.1 (RD = -1)",
    "D22.1 (RD = +1)",
    "D23.1 (RD = -1)",
    "D23.1 (RD = +1)",
    "D24.1 (RD = -1)",
    "D24.1 (RD = +1)",
    "D25.1 (RD = -1)",
    "D25.1 (RD = +1)",
    "D26.1 (RD = -1)",
    "D26.1 (RD = +1)",
    "D27.1 (RD = -1)",
    "D27.1 (RD = +1)",
    "D28.1 (RD = -1)",
    "D28.1 (RD = +1)",
    "D29.1 (RD = -1)",
    "D29.1 (RD = +1)",
    "D30.1 (RD = -1)",
    "D30.1 (RD = +1)",
    "D31.1 (RD = -1)",
    "D31.1 (RD = +1)",
    "D00.2 (RD = -1)",
    "D00.2 (RD = +1)",
    "D01.2 (RD = -1)",
    "D01.2 (RD = +1)",
    "D02.2 (RD = -1)",
    "D02.2 (RD = +1)",
    "D03.2 (RD = -1)",
    "D03.2 (RD = +1)",
    "D04.2 (RD = -1)",
    "D04.2 (RD = +1)",
    "D05.2 (RD = -1)",
    "D05.2 (RD = +1)",
    "D06.2 (RD = -1)",
    "D06.2 (RD = +1)",
    "D07.2 (RD = -1)",
    "D07.2 (RD = +1)",
    "D08.2 (RD = -1)",
    "D08.2 (RD = +1)",
    "D09.2 (RD = -1)",
    "D09.2 (RD = +1)",
    "D10.2 (RD = -1)",
    "D10.2 (RD = +1)",
    "D11.2 (RD = -1)",
    "D11.2 (RD = +1)",
    "D12.2 (RD = -1)",
    "D12.2 (RD = +1)",
    "D13.2 (RD = -1)",
    "D13.2 (RD = +1)",
    "D14.2 (RD = -1)",
    "D14.2 (RD = +1)",
    "D15.2 (RD = -1)",
    "D15.2 (RD = +1)",
    "D16.2 (RD = -1)",
    "D16.2 (RD = +1)",
    "D17.2 (RD = -1)",
    "D17.2 (RD = +1)",
    "D18.2 (RD = -1)",
    "D18.2 (RD = +1)",
    "D19.2 (RD = -1)",
    "D19.2 (RD = +1)",
    "D20.2 (RD = -1)",
    "D20.2 (RD = +1)",
    "D21.2 (RD = -1)",
    "D21.2 (RD = +1)",
    "D22.2 (RD = -1)",
    "D22.2 (RD = +1)",
    "D23.2 (RD = -1)",
    "D23.2 (RD = +1)",
    "D24.2 (RD = -1)",
    "D24.2 (RD = +1)",
    "D25.2 (RD = -1)",
    "D25.2 (RD = +1)",
    "D26.2 (RD = -1)",
    "D26.2 (RD = +1)",
    "D27.2 (RD = -1)",
    "D27.2 (RD = +1)",
    "D28.2 (RD = -1)",
    "D28.2 (RD = +1)",
    "D29.2 (RD = -1)",
    "D29.2 (RD = +1)",
    "D30.2 (RD = -1)",
    "D30.2 (RD = +1)",
    "D31.2 (RD = -1)",
    "D31.2 (RD = +1)",
    "D00.3 (RD = -1)",
    "D00.3 (RD = +1)",
    "D01.3 (RD = -1)",
    "D01.3 (RD = +1)",
    "D02.3 (RD = -1)",
    "D02.3 (RD = +1)",
    "D03.3 (RD = -1)",
    "D03.3 (RD = +1)",
    "D04.3 (RD = -1)",
    "D04.3 (RD = +1)",
    "D05.3 (RD = -1)",
    "D05.3 (RD = +1)",
    "D06.3 (RD = -1)",
    "D06.3 (RD = +1)",
    "D07.3 (RD = -1)",
    "D07.3 (RD = +1)",
    "D08.3 (RD = -1)",
    "D08.3 (RD = +1)",
    "D09.3 (RD = -1)",
    "D09.3 (RD = +1)",
    "D10.3 (RD = -1)",
    "D10.3 (RD = +1)",
    "D11.3 (RD = -1)",
    "D11.3 (RD = +1)",
    "D12.3 (RD = -1)",
    "D12.3 (RD = +1)",
    "D13.3 (RD = -1)",
    "D13.3 (RD = +1)",
    "D14.3 (RD = -1)",
    "D14.3 (RD = +1)",
    "D15.3 (RD = -1)",
    "D15.3 (RD = +1)",
    "D16.3 (RD = -1)",
    "D16.3 (RD = +1)",
    "D17.3 (RD = -1)",
    "D17.3 (RD = +1)",
    "D18.3 (RD = -1)",
    "D18.3 (RD = +1)",
    "D19.3 (RD = -1)",
    "D19.3 (RD = +1)",
    "D20.3 (RD = -1)",
    "D20.3 (RD = +1)",
    "D21.3 (RD = -1)",
    "D21.3 (RD = +1)",
    "D22.3 (RD = -1)",
    "D22.3 (RD = +1)",
    "D23.3 (RD = -1)",
    "D23.3 (RD = +1)",
    "D24.3 (RD = -1)",
    "D24.3 (RD = +1)",
    "D25.3 (RD = -1)",
    "D25.3 (RD = +1)",
    "D26.3 (RD = -1)",
    "D26.3 (RD = +1)",
    "D27.3 (RD = -1)",
    "D27.3 (RD = +1)",
    "D28.3 (RD = -1)",
    "D28.3 (RD = +1)",
    "D29.3 (RD = -1)",
    "D29.3 (RD = +1)",
    "D30.3 (RD = -1)",
    "D30.3 (RD = +1)",
    "D31.3 (RD = -1)",
    "D31.3 (RD = +1)",
    "D00.4 (RD = -1)",
    "D00.4 (RD = +1)",
    "D01.4 (RD = -1)",
    "D01.4 (RD = +1)",
    "D02.4 (RD = -1)",
    "D02.4 (RD = +1)",
    "D03.4 (RD = -1)",
    "D03.4 (RD = +1)",
    "D04.4 (RD = -1)",
    "D04.4 (RD = +1)",
    "D05.4 (RD = -1)",
    "D05.4 (RD = +1)",
    "D06.4 (RD = -1)",
    "D06.4 (RD = +1)",
    "D07.4 (RD = -1)",
    "D07.4 (RD = +1)",
    "D08.4 (RD = -1)",
    "D08.4 (RD = +1)",
    "D09.4 (RD = -1)",
    "D09.4 (RD = +1)",
    "D10.4 (RD = -1)",
    "D10.4 (RD = +1)",
    "D11.4 (RD = -1)",
    "D11.4 (RD = +1)",
    "D12.4 (RD = -1)",
    "D12.4 (RD = +1)",
    "D13.4 (RD = -1)",
    "D13.4 (RD = +1)",
    "D14.4 (RD = -1)",
    "D14.4 (RD = +1)",
    "D15.4 (RD = -1)",
    "D15.4 (RD = +1)",
    "D16.4 (RD = -1)",
    "D16.4 (RD = +1)",
    "D17.4 (RD = -1)",
    "D17.4 (RD = +1)",
    "D18.4 (RD = -1)",
    "D18.4 (RD = +1)",
    "D19.4 (RD = -1)",
    "D19.4 (RD = +1)",
    "D20.4 (RD = -1)",
    "D20.4 (RD = +1)",
    "D21.4 (RD = -1)",
    "D21.4 (RD = +1)",
    "D22.4 (RD = -1)",
    "D22.4 (RD = +1)",
    "D23.4 (RD = -1)",
    "D23.4 (RD = +1)",
    "D24.4 (RD = -1)",
    "D24.4 (RD = +1)",
    "D25.4 (RD = -1)",
    "D25.4 (RD = +1)",
    "D26.4 (RD = -1)",
    "D26.4 (RD = +1)",
    "D27.4 (RD = -1)",
    "D27.4 (RD = +1)",
    "D28.4 (RD = -1)",
    "D28.4 (RD = +1)",
    "D29.4 (RD = -1)",
    "D29.4 (RD = +1)",
    "D30.4 (RD = -1)",
    "D30.4 (RD = +1)",
    "D31.4 (RD = -1)",
    "D31.4 (RD = +1)",
    "D00.5 (RD = -1)",
    "D00.5 (RD = +1)",
    "D01.5 (RD = -1)",
    "D01.5 (RD = +1)",
    "D02.5 (RD = -1)",
    "D02.5 (RD = +1)",
    "D03.5 (RD = -1)",
    "D03.5 (RD = +1)",
    "D04.5 (RD = -1)",
    "D04.5 (RD = +1)",
    "D05.5 (RD = -1)",
    "D05.5 (RD = +1)",
    "D06.5 (RD = -1)",
    "D06.5 (RD = +1)",
    "D07.5 (RD = -1)",
    "D07.5 (RD = +1)",
    "D08.5 (RD = -1)",
    "D08.5 (RD = +1)",
    "D09.5 (RD = -1)",
    "D09.5 (RD = +1)",
    "D10.5 (RD = -1)",
    "D10.5 (RD = +1)",
    "D11.5 (RD = -1)",
    "D11.5 (RD = +1)",
    "D12.5 (RD = -1)",
    "D12.5 (RD = +1)",
    "D13.5 (RD = -1)",
    "D13.5 (RD = +1)",
    "D14.5 (RD = -1)",
    "D14.5 (RD = +1)",
    "D15.5 (RD = -1)",
    "D15.5 (RD = +1)",
    "D16.5 (RD = -1)",
    "D16.5 (RD = +1)",
    "D17.5 (RD = -1)",
    "D17.5 (RD = +1)",
    "D18.5 (RD = -1)",
    "D18.5 (RD = +1)",
    "D19.5 (RD = -1)",
    "D19.5 (RD = +1)",
    "D20.5 (RD = -1)",
    "D20.5 (RD = +1)",
    "D21.5 (RD = -1)",
    "D21.5 (RD = +1)",
    "D22.5 (RD = -1)",
    "D22.5 (RD = +1)",
    "D23.5 (RD = -1)",
    "D23.5 (RD = +1)",
    "D24.5 (RD = -1)",
    "D24.5 (RD = +1)",
    "D25.5 (RD = -1)",
    "D25.5 (RD = +1)",
    "D26.5 (RD = -1)",
    "D26.5 (RD = +1)",
    "D27.5 (RD = -1)",
    "D27.5 (RD = +1)",
    "D28.5 (RD = -1)",
    "D28.5 (RD = +1)",
    "D29.5 (RD = -1)",
    "D29.5 (RD = +1)",
    "D30.5 (RD = -1)",
    "D30.5 (RD = +1)",
    "D31.5 (RD = -1)",
    "D31.5 (RD = +1)",
    "D00.6 (RD = -1)",
    "D00.6 (RD = +1)",
    "D01.6 (RD = -1)",
    "D01.6 (RD = +1)",
    "D02.6 (RD = -1)",
    "D02.6 (RD = +1)",
    "D03.6 (RD = -1)",
    "D03.6 (RD = +1)",
    "D04.6 (RD = -1)",
    "D04.6 (RD = +1)",
    "D05.6 (RD = -1)",
    "D05.6 (RD = +1)",
    "D06.6 (RD = -1)",
    "D06.6 (RD = +1)",
    "D07.6 (RD = -1)",
    "D07.6 (RD = +1)",
    "D08.6 (RD = -1)",
    "D08.6 (RD = +1)",
    "D09.6 (RD = -1)",
    "D09.6 (RD = +1)",
    "D10.6 (RD = -1)",
    "D10.6 (RD = +1)",
    "D11.6 (RD = -1)",
    "D11.6 (RD = +1)",
    "D12.6 (RD = -1)",
    "D12.6 (RD = +1)",
    "D13.6 (RD = -1)",
    "D13.6 (RD = +1)",
    "D14.6 (RD = -1)",
    "D14.6 (RD = +1)",
    "D15.6 (RD = -1)",
    "D15.6 (RD = +1)",
    "D16.6 (RD = -1)",
    "D16.6 (RD = +1)",
    "D17.6 (RD = -1)",
    "D17.6 (RD = +1)",
    "D18.6 (RD = -1)",
    "D18.6 (RD = +1)",
    "D19.6 (RD = -1)",
    "D19.6 (RD = +1)",
    "D20.6 (RD = -1)",
    "D20.6 (RD = +1)",
    "D21.6 (RD = -1)",
    "D21.6 (RD = +1)",
    "D22.6 (RD = -1)",
    "D22.6 (RD = +1)",
    "D23.6 (RD = -1)",
    "D23.6 (RD = +1)",
    "D24.6 (RD = -1)",
    "D24.6 (RD = +1)",
    "D25.6 (RD = -1)",
    "D25.6 (RD = +1)",
    "D26.6 (RD = -1)",
    "D26.6 (RD = +1)",
    "D27.6 (RD = -1)",
    "D27.6 (RD = +1)",
    "D28.6 (RD = -1)",
    "D28.6 (RD = +1)",
    "D29.6 (RD = -1)",
    "D29.6 (RD = +1)",
    "D30.6 (RD = -1)",
    "D30.6 (RD = +1)",
    "D31.6 (RD = -1)",
    "D31.6 (RD = +1)",
    "D00.7 (RD = -1)",
    "D00.7 (RD = +1)",
    "D01.7 (RD = -1)",
    "D01.7 (RD = +1)",
    "D02.7 (RD = -1)",
    "D02.7 (RD = +1)",
    "D03.7 (RD = -1)",
    "D03.7 (RD = +1)",
    "D04.7 (RD = -1)",
    "D04.7 (RD = +1)",
    "D05.7 (RD = -1)",
    "D05.7 (RD = +1)",
    "D06.7 (RD = -1)",
    "D06.7 (RD = +1)",
    "D07.7 (RD = -1)",
    "D07.7 (RD = +1)",
    "D08.7 (RD = -1)",
    "D08.7 (RD = +1)",
    "D09.7 (RD = -1)",
    "D09.7 (RD = +1)",
    "D10.7 (RD = -1)",
    "D10.7 (RD = +1)",
    "D11.7 (RD = -1)",
    "D11.7 (RD = +1)",
    "D12.7 (RD = -1)",
    "D12.7 (RD = +1)",
    "D13.7 (RD = -1)",
    "D13.7 (RD = +1)",
    "D14.7 (RD = -1)",
    "D14.7 (RD = +1)",
    "D15.7 (RD = -1)",
    "D15.7 (RD = +1)",
    "D16.7 (RD = -1)",
    "D16.7 (RD = +1)",
    "D17.7 (RD = -1)",
    "D17.7 (RD = +1)",
    "D18.7 (RD = -1)",
    "D18.7 (RD = +1)",
    "D19.7 (RD = -1)",
    "D19.7 (RD = +1)",
    "D20.7 (RD = -1)",
    "D20.7 (RD = +1)",
    "D21.7 (RD = -1)",
    "D21.7 (RD = +1)",
    "D22.7 (RD = -1)",
    "D22.7 (RD = +1)",
    "D23.7 (RD = -1)",
    "D23.7 (RD = +1)",
    "D24.7 (RD = -1)",
    "D24.7 (RD = +1)",
    "D25.7 (RD = -1)",
    "D25.7 (RD = +1)",
    "D26.7 (RD = -1)",
    "D26.7 (RD = +1)",
    "D27.7 (RD = -1)",
    "D27.7 (RD = +1)",
    "D28.7 (RD = -1)",
    "D28.7 (RD = +1)",
    "D29.7 (RD = -1)",
    "D29.7 (RD = +1)",
    "D30.7 (RD = -1)",
    "D30.7 (RD = +1)",
    "D31.7 (RD = -1)",
    "D31.7 (RD = +1)",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "K28.0 (RD = -1)",
    "K28.0 (RD = +1)",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "K28.1 (RD = -1)",
    "K28.1 (RD = +1)",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "K28.2 (RD = -1)",
    "K28.2 (RD = +1)",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "K28.3 (RD = -1)",
    "K28.3 (RD = +1)",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "K28.4 (RD = -1)",
    "K28.4 (RD = +1)",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "K28.5 (RD = -1)",
    "K28.5 (RD = +1)",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "K28.6 (RD = -1)",
    "K28.6 (RD = +1)",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "K23.7 (RD = -1)",
    "K23.7 (RD = +1)",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "K27.7 (RD = -1)",
    "K27.7 (RD = +1)",
    "K28.7 (RD = -1)",
    "K28.7 (RD = +1)",
    "K29.7 (RD = -1)",
    "K29.7 (RD = +1)",
    "K30.7 (RD = -1)",
    "K30.7 (RD = +1)",
    "?",
    "?"
  };

  logic [1+1+1+2+8+10+2-1:0] dec_table [2048] = '{
    //DV   WRONG K     RDF    octet        code            RDE
    //24   23    22    21:20  19:12        11:2            1:0
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0000000000, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0000000001, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0000000010, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0000000011, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0000000100, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0000000101, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0000000110, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0000000111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0000001000, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0000001001, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0000001010, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0000001011, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0000001100, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0000001101, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0000001110, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0000001111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0000010000, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0000010001, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0000010010, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0000010011, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0000010100, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0000010101, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0000010110, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0000010111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0000011000, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0000011001, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0000011010, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0000011011, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0000011100, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0000011101, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0000011110, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0000011111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0000100000, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0000100001, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0000100010, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0000100011, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0000100100, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0000100101, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0000100110, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0000100111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0000101000, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0000101001, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0000101010, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0000101011, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0000101100, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0000101101, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0000101110, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0000101111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0000110000, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0000110001, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0000110010, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0000110011, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0000110100, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0000110101, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0000110110, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0000110111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0000111000, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0000111001, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0000111010, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0000111011, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0000111100, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0000111101, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0000111110, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0000111111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0001000000, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0001000001, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0001000010, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0001000011, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0001000100, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0001000101, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0001000110, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0001000111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0001001000, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0001001001, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0001001010, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0001001011, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0001001100, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0001001101, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0001001110, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0001001111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0001010000, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0001010001, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0001010010, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0001010011, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0001010100, 2'bxx}, // ?
    {1'b1, 1'b0, 1'b0, 2'b11, 8'b01010111, 10'b0001010101, 2'b11}, // D23.2 (RD = +1) WRONG RDF
    {1'b1, 1'b0, 1'b0, 2'b11, 8'b11010111, 10'b0001010110, 2'b11}, // D23.6 (RD = +1) WRONG RDF
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0001010111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0001011000, 2'bxx}, // ?
    {1'b1, 1'b0, 1'b0, 2'b11, 8'b00110111, 10'b0001011001, 2'b11}, // D23.1 (RD = +1) WRONG RDF
    {1'b1, 1'b0, 1'b0, 2'b11, 8'b10110111, 10'b0001011010, 2'b11}, // D23.5 (RD = +1) WRONG RDF
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0001011011, 2'bxx}, // ?
    {1'b1, 1'b0, 1'b0, 2'b11, 8'b01110111, 10'b0001011100, 2'b11}, // D23.3 (RD = +1) WRONG RDF
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0001011101, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0001011110, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0001011111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0001100000, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0001100001, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0001100010, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0001100011, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0001100100, 2'bxx}, // ?
    {1'b1, 1'b0, 1'b0, 2'b11, 8'b01001000, 10'b0001100101, 2'b11}, // D08.2 (RD = +1) WRONG RDF
    {1'b1, 1'b0, 1'b0, 2'b11, 8'b11001000, 10'b0001100110, 2'b11}, // D08.6 (RD = +1) WRONG RDF
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0001100111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0001101000, 2'bxx}, // ?
    {1'b1, 1'b0, 1'b0, 2'b11, 8'b00101000, 10'b0001101001, 2'b11}, // D08.1 (RD = +1) WRONG RDF
    {1'b1, 1'b0, 1'b0, 2'b11, 8'b10101000, 10'b0001101010, 2'b11}, // D08.5 (RD = +1) WRONG RDF
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0001101011, 2'bxx}, // ?
    {1'b1, 1'b0, 1'b0, 2'b11, 8'b01101000, 10'b0001101100, 2'b11}, // D08.3 (RD = +1) WRONG RDF
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0001101101, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0001101110, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0001101111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0001110000, 2'bxx}, // ?
    {1'b1, 1'b0, 1'b0, 2'b11, 8'b11100111, 10'b0001110001, 2'b11}, // D07.7 (RD = +1) WRONG RDF
    {1'b1, 1'b0, 1'b0, 2'b11, 8'b10000111, 10'b0001110010, 2'b11}, // D07.4 (RD = +1) WRONG RDF
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0001110011, 2'bxx}, // ?
    {1'b1, 1'b0, 1'b0, 2'b11, 8'b00000111, 10'b0001110100, 2'b11}, // D07.0 (RD = +1) WRONG RDF
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0001110101, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0001110110, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0001110111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0001111000, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0001111001, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0001111010, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0001111011, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0001111100, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0001111101, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0001111110, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0001111111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0010000000, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0010000001, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0010000010, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0010000011, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0010000100, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0010000101, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0010000110, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0010000111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0010001000, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0010001001, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0010001010, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0010001011, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0010001100, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0010001101, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0010001110, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0010001111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0010010000, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0010010001, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0010010010, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0010010011, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0010010100, 2'bxx}, // ?
    {1'b1, 1'b0, 1'b0, 2'b11, 8'b01011011, 10'b0010010101, 2'b11}, // D27.2 (RD = +1) WRONG RDF
    {1'b1, 1'b0, 1'b0, 2'b11, 8'b11011011, 10'b0010010110, 2'b11}, // D27.6 (RD = +1) WRONG RDF
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0010010111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0010011000, 2'bxx}, // ?
    {1'b1, 1'b0, 1'b0, 2'b11, 8'b00111011, 10'b0010011001, 2'b11}, // D27.1 (RD = +1) WRONG RDF
    {1'b1, 1'b0, 1'b0, 2'b11, 8'b10111011, 10'b0010011010, 2'b11}, // D27.5 (RD = +1) WRONG RDF
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0010011011, 2'bxx}, // ?
    {1'b1, 1'b0, 1'b0, 2'b11, 8'b01111011, 10'b0010011100, 2'b11}, // D27.3 (RD = +1) WRONG RDF
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0010011101, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0010011110, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0010011111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0010100000, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0010100001, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0010100010, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0010100011, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0010100100, 2'bxx}, // ?
    {1'b1, 1'b0, 1'b0, 2'b11, 8'b01000100, 10'b0010100101, 2'b11}, // D04.2 (RD = +1) WRONG RDF
    {1'b1, 1'b0, 1'b0, 2'b11, 8'b11000100, 10'b0010100110, 2'b11}, // D04.6 (RD = +1) WRONG RDF
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0010100111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0010101000, 2'bxx}, // ?
    {1'b1, 1'b0, 1'b0, 2'b11, 8'b00100100, 10'b0010101001, 2'b11}, // D04.1 (RD = +1) WRONG RDF
    {1'b1, 1'b0, 1'b0, 2'b11, 8'b10100100, 10'b0010101010, 2'b11}, // D04.5 (RD = +1) WRONG RDF
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0010101011, 2'bxx}, // ?
    {1'b1, 1'b0, 1'b0, 2'b11, 8'b01100100, 10'b0010101100, 2'b11}, // D04.3 (RD = +1) WRONG RDF
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0010101101, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0010101110, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0010101111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0010110000, 2'bxx}, // ?
    {1'b1, 1'b0, 1'b0, 2'b11, 8'b11110100, 10'b0010110001, 2'b11}, // D20.7 (RD = +1) WRONG RDF
    {1'b1, 1'b0, 1'b0, 2'b11, 8'b10010100, 10'b0010110010, 2'b11}, // D20.4 (RD = +1) WRONG RDF
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0010110011, 2'bxx}, // ?
    {1'b1, 1'b0, 1'b0, 2'b11, 8'b00010100, 10'b0010110100, 2'b11}, // D20.0 (RD = +1) WRONG RDF
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b01010100, 10'b0010110101, 2'b11}, // D20.2 (RD = -1)
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b11010100, 10'b0010110110, 2'b11}, // D20.6 (RD = -1)
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b11110100, 10'b0010110111, 2'b01}, // D20.7 (RD = -1)
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0010111000, 2'bxx}, // ?
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b00110100, 10'b0010111001, 2'b11}, // D20.1 (RD = -1)
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b10110100, 10'b0010111010, 2'b11}, // D20.5 (RD = -1)
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b00010100, 10'b0010111011, 2'b01}, // D20.0 (RD = -1)
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b01110100, 10'b0010111100, 2'b11}, // D20.3 (RD = -1)
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b10010100, 10'b0010111101, 2'b01}, // D20.4 (RD = -1)
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0010111110, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0010111111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0011000000, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0011000001, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0011000010, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0011000011, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0011000100, 2'bxx}, // ?
    {1'b1, 1'b0, 1'b0, 2'b11, 8'b01011000, 10'b0011000101, 2'b11}, // D24.2 (RD = +1) WRONG RDF
    {1'b1, 1'b0, 1'b0, 2'b11, 8'b11011000, 10'b0011000110, 2'b11}, // D24.6 (RD = +1) WRONG RDF
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0011000111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0011001000, 2'bxx}, // ?
    {1'b1, 1'b0, 1'b0, 2'b11, 8'b00111000, 10'b0011001001, 2'b11}, // D24.1 (RD = +1) WRONG RDF
    {1'b1, 1'b0, 1'b0, 2'b11, 8'b10111000, 10'b0011001010, 2'b11}, // D24.5 (RD = +1) WRONG RDF
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0011001011, 2'bxx}, // ?
    {1'b1, 1'b0, 1'b0, 2'b11, 8'b01111000, 10'b0011001100, 2'b11}, // D24.3 (RD = +1) WRONG RDF
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0011001101, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0011001110, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0011001111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0011010000, 2'bxx}, // ?
    {1'b1, 1'b0, 1'b0, 2'b11, 8'b11101100, 10'b0011010001, 2'b11}, // D12.7 (RD = +1) WRONG RDF
    {1'b1, 1'b0, 1'b0, 2'b11, 8'b10001100, 10'b0011010010, 2'b11}, // D12.4 (RD = +1) WRONG RDF
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0011010011, 2'bxx}, // ?
    {1'b1, 1'b0, 1'b0, 2'b11, 8'b00001100, 10'b0011010100, 2'b11}, // D12.0 (RD = +1) WRONG RDF
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b01001100, 10'b0011010101, 2'b11}, // D12.2 (RD = -1)
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b11001100, 10'b0011010110, 2'b11}, // D12.6 (RD = -1)
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0011010111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0011011000, 2'bxx}, // ?
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b00101100, 10'b0011011001, 2'b11}, // D12.1 (RD = -1)
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b10101100, 10'b0011011010, 2'b11}, // D12.5 (RD = -1)
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b00001100, 10'b0011011011, 2'b01}, // D12.0 (RD = -1)
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b01101100, 10'b0011011100, 2'b11}, // D12.3 (RD = -1)
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b10001100, 10'b0011011101, 2'b01}, // D12.4 (RD = -1)
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b11101100, 10'b0011011110, 2'b01}, // D12.7 (RD = -1)
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0011011111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0011100000, 2'bxx}, // ?
    {1'b1, 1'b0, 1'b0, 2'b11, 8'b11111100, 10'b0011100001, 2'b11}, // D28.7 (RD = +1) WRONG RDF
    {1'b1, 1'b0, 1'b0, 2'b11, 8'b10011100, 10'b0011100010, 2'b11}, // D28.4 (RD = +1) WRONG RDF
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0011100011, 2'bxx}, // ?
    {1'b1, 1'b0, 1'b0, 2'b11, 8'b00011100, 10'b0011100100, 2'b11}, // D28.0 (RD = +1) WRONG RDF
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b01011100, 10'b0011100101, 2'b11}, // D28.2 (RD = -1)
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b11011100, 10'b0011100110, 2'b11}, // D28.6 (RD = -1)
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0011100111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0011101000, 2'bxx}, // ?
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b00111100, 10'b0011101001, 2'b11}, // D28.1 (RD = -1)
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b10111100, 10'b0011101010, 2'b11}, // D28.5 (RD = -1)
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b00011100, 10'b0011101011, 2'b01}, // D28.0 (RD = -1)
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b01111100, 10'b0011101100, 2'b11}, // D28.3 (RD = -1)
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b10011100, 10'b0011101101, 2'b01}, // D28.4 (RD = -1)
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b11111100, 10'b0011101110, 2'b01}, // D28.7 (RD = -1)
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0011101111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0011110000, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0011110001, 2'bxx}, // ?
    {1'b0, 1'b0, 1'b1, 2'b11, 8'b10011100, 10'b0011110010, 2'b11}, // K28.4 (RD = -1)
    {1'b0, 1'b0, 1'b1, 2'b11, 8'b01111100, 10'b0011110011, 2'b01}, // K28.3 (RD = -1)
    {1'b0, 1'b0, 1'b1, 2'b11, 8'b00011100, 10'b0011110100, 2'b11}, // K28.0 (RD = -1)
    {1'b0, 1'b0, 1'b1, 2'b11, 8'b01011100, 10'b0011110101, 2'b01}, // K28.2 (RD = -1)
    {1'b0, 1'b0, 1'b1, 2'b11, 8'b11011100, 10'b0011110110, 2'b01}, // K28.6 (RD = -1)
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0011110111, 2'bxx}, // ?
    {1'b0, 1'b0, 1'b1, 2'b11, 8'b11111100, 10'b0011111000, 2'b11}, // K28.7 (RD = -1)
    {1'b0, 1'b0, 1'b1, 2'b11, 8'b00111100, 10'b0011111001, 2'b01}, // K28.1 (RD = -1)
    {1'b0, 1'b0, 1'b1, 2'b11, 8'b10111100, 10'b0011111010, 2'b01}, // K28.5 (RD = -1)
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0011111011, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0011111100, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0011111101, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0011111110, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0011111111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0100000000, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0100000001, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0100000010, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0100000011, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0100000100, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0100000101, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0100000110, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0100000111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0100001000, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0100001001, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0100001010, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0100001011, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0100001100, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0100001101, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0100001110, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0100001111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0100010000, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0100010001, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0100010010, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0100010011, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0100010100, 2'bxx}, // ?
    {1'b1, 1'b0, 1'b0, 2'b11, 8'b01011101, 10'b0100010101, 2'b11}, // D29.2 (RD = +1) WRONG RDF
    {1'b1, 1'b0, 1'b0, 2'b11, 8'b11011101, 10'b0100010110, 2'b11}, // D29.6 (RD = +1) WRONG RDF
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0100010111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0100011000, 2'bxx}, // ?
    {1'b1, 1'b0, 1'b0, 2'b11, 8'b00111101, 10'b0100011001, 2'b11}, // D29.1 (RD = +1) WRONG RDF
    {1'b1, 1'b0, 1'b0, 2'b11, 8'b10111101, 10'b0100011010, 2'b11}, // D29.5 (RD = +1) WRONG RDF
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0100011011, 2'bxx}, // ?
    {1'b1, 1'b0, 1'b0, 2'b11, 8'b01111101, 10'b0100011100, 2'b11}, // D29.3 (RD = +1) WRONG RDF
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0100011101, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0100011110, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0100011111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0100100000, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0100100001, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0100100010, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0100100011, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0100100100, 2'bxx}, // ?
    {1'b1, 1'b0, 1'b0, 2'b11, 8'b01000010, 10'b0100100101, 2'b11}, // D02.2 (RD = +1) WRONG RDF
    {1'b1, 1'b0, 1'b0, 2'b11, 8'b11000010, 10'b0100100110, 2'b11}, // D02.6 (RD = +1) WRONG RDF
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0100100111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0100101000, 2'bxx}, // ?
    {1'b1, 1'b0, 1'b0, 2'b11, 8'b00100010, 10'b0100101001, 2'b11}, // D02.1 (RD = +1) WRONG RDF
    {1'b1, 1'b0, 1'b0, 2'b11, 8'b10100010, 10'b0100101010, 2'b11}, // D02.5 (RD = +1) WRONG RDF
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0100101011, 2'bxx}, // ?
    {1'b1, 1'b0, 1'b0, 2'b11, 8'b01100010, 10'b0100101100, 2'b11}, // D02.3 (RD = +1) WRONG RDF
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0100101101, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0100101110, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0100101111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0100110000, 2'bxx}, // ?
    {1'b1, 1'b0, 1'b0, 2'b11, 8'b11110010, 10'b0100110001, 2'b11}, // D18.7 (RD = +1) WRONG RDF
    {1'b1, 1'b0, 1'b0, 2'b11, 8'b10010010, 10'b0100110010, 2'b11}, // D18.4 (RD = +1) WRONG RDF
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0100110011, 2'bxx}, // ?
    {1'b1, 1'b0, 1'b0, 2'b11, 8'b00010010, 10'b0100110100, 2'b11}, // D18.0 (RD = +1) WRONG RDF
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b01010010, 10'b0100110101, 2'b11}, // D18.2 (RD = -1)
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b11010010, 10'b0100110110, 2'b11}, // D18.6 (RD = -1)
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b11110010, 10'b0100110111, 2'b01}, // D18.7 (RD = -1)
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0100111000, 2'bxx}, // ?
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b00110010, 10'b0100111001, 2'b11}, // D18.1 (RD = -1)
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b10110010, 10'b0100111010, 2'b11}, // D18.5 (RD = -1)
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b00010010, 10'b0100111011, 2'b01}, // D18.0 (RD = -1)
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b01110010, 10'b0100111100, 2'b11}, // D18.3 (RD = -1)
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b10010010, 10'b0100111101, 2'b01}, // D18.4 (RD = -1)
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0100111110, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0100111111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0101000000, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0101000001, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0101000010, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0101000011, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0101000100, 2'bxx}, // ?
    {1'b1, 1'b0, 1'b0, 2'b11, 8'b01011111, 10'b0101000101, 2'b11}, // D31.2 (RD = +1) WRONG RDF
    {1'b1, 1'b0, 1'b0, 2'b11, 8'b11011111, 10'b0101000110, 2'b11}, // D31.6 (RD = +1) WRONG RDF
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0101000111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0101001000, 2'bxx}, // ?
    {1'b1, 1'b0, 1'b0, 2'b11, 8'b00111111, 10'b0101001001, 2'b11}, // D31.1 (RD = +1) WRONG RDF
    {1'b1, 1'b0, 1'b0, 2'b11, 8'b10111111, 10'b0101001010, 2'b11}, // D31.5 (RD = +1) WRONG RDF
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0101001011, 2'bxx}, // ?
    {1'b1, 1'b0, 1'b0, 2'b11, 8'b01111111, 10'b0101001100, 2'b11}, // D31.3 (RD = +1) WRONG RDF
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0101001101, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0101001110, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0101001111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0101010000, 2'bxx}, // ?
    {1'b1, 1'b0, 1'b0, 2'b11, 8'b11101010, 10'b0101010001, 2'b11}, // D10.7 (RD = +1) WRONG RDF
    {1'b1, 1'b0, 1'b0, 2'b11, 8'b10001010, 10'b0101010010, 2'b11}, // D10.4 (RD = +1) WRONG RDF
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0101010011, 2'bxx}, // ?
    {1'b1, 1'b0, 1'b0, 2'b11, 8'b00001010, 10'b0101010100, 2'b11}, // D10.0 (RD = +1) WRONG RDF
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b01001010, 10'b0101010101, 2'b11}, // D10.2 (RD = -1)
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b11001010, 10'b0101010110, 2'b11}, // D10.6 (RD = -1)
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0101010111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0101011000, 2'bxx}, // ?
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b00101010, 10'b0101011001, 2'b11}, // D10.1 (RD = -1)
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b10101010, 10'b0101011010, 2'b11}, // D10.5 (RD = -1)
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b00001010, 10'b0101011011, 2'b01}, // D10.0 (RD = -1)
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b01101010, 10'b0101011100, 2'b11}, // D10.3 (RD = -1)
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b10001010, 10'b0101011101, 2'b01}, // D10.4 (RD = -1)
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b11101010, 10'b0101011110, 2'b01}, // D10.7 (RD = -1)
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0101011111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0101100000, 2'bxx}, // ?
    {1'b1, 1'b0, 1'b0, 2'b11, 8'b11111010, 10'b0101100001, 2'b11}, // D26.7 (RD = +1) WRONG RDF
    {1'b1, 1'b0, 1'b0, 2'b11, 8'b10011010, 10'b0101100010, 2'b11}, // D26.4 (RD = +1) WRONG RDF
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0101100011, 2'bxx}, // ?
    {1'b1, 1'b0, 1'b0, 2'b11, 8'b00011010, 10'b0101100100, 2'b11}, // D26.0 (RD = +1) WRONG RDF
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b01011010, 10'b0101100101, 2'b11}, // D26.2 (RD = -1)
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b11011010, 10'b0101100110, 2'b11}, // D26.6 (RD = -1)
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0101100111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0101101000, 2'bxx}, // ?
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b00111010, 10'b0101101001, 2'b11}, // D26.1 (RD = -1)
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b10111010, 10'b0101101010, 2'b11}, // D26.5 (RD = -1)
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b00011010, 10'b0101101011, 2'b01}, // D26.0 (RD = -1)
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b01111010, 10'b0101101100, 2'b11}, // D26.3 (RD = -1)
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b10011010, 10'b0101101101, 2'b01}, // D26.4 (RD = -1)
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b11111010, 10'b0101101110, 2'b01}, // D26.7 (RD = -1)
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0101101111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0101110000, 2'bxx}, // ?
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b11101111, 10'b0101110001, 2'b11}, // D15.7 (RD = -1)
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b10001111, 10'b0101110010, 2'b11}, // D15.4 (RD = -1)
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b01101111, 10'b0101110011, 2'b01}, // D15.3 (RD = -1)
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b00001111, 10'b0101110100, 2'b11}, // D15.0 (RD = -1)
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b01001111, 10'b0101110101, 2'b01}, // D15.2 (RD = -1)
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b11001111, 10'b0101110110, 2'b01}, // D15.6 (RD = -1)
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0101110111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0101111000, 2'bxx}, // ?
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b00101111, 10'b0101111001, 2'b01}, // D15.1 (RD = -1)
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b10101111, 10'b0101111010, 2'b01}, // D15.5 (RD = -1)
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0101111011, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0101111100, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0101111101, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0101111110, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0101111111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0110000000, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0110000001, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0110000010, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0110000011, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0110000100, 2'bxx}, // ?
    {1'b1, 1'b0, 1'b0, 2'b11, 8'b01000000, 10'b0110000101, 2'b11}, // D00.2 (RD = +1) WRONG RDF
    {1'b1, 1'b0, 1'b0, 2'b11, 8'b11000000, 10'b0110000110, 2'b11}, // D00.6 (RD = +1) WRONG RDF
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0110000111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0110001000, 2'bxx}, // ?
    {1'b1, 1'b0, 1'b0, 2'b11, 8'b00100000, 10'b0110001001, 2'b11}, // D00.1 (RD = +1) WRONG RDF
    {1'b1, 1'b0, 1'b0, 2'b11, 8'b10100000, 10'b0110001010, 2'b11}, // D00.5 (RD = +1) WRONG RDF
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0110001011, 2'bxx}, // ?
    {1'b1, 1'b0, 1'b0, 2'b11, 8'b01100000, 10'b0110001100, 2'b11}, // D00.3 (RD = +1) WRONG RDF
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0110001101, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0110001110, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0110001111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0110010000, 2'bxx}, // ?
    {1'b1, 1'b0, 1'b0, 2'b11, 8'b11100110, 10'b0110010001, 2'b11}, // D06.7 (RD = +1) WRONG RDF
    {1'b1, 1'b0, 1'b0, 2'b11, 8'b10000110, 10'b0110010010, 2'b11}, // D06.4 (RD = +1) WRONG RDF
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0110010011, 2'bxx}, // ?
    {1'b1, 1'b0, 1'b0, 2'b11, 8'b00000110, 10'b0110010100, 2'b11}, // D06.0 (RD = +1) WRONG RDF
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b01000110, 10'b0110010101, 2'b11}, // D06.2 (RD = -1)
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b11000110, 10'b0110010110, 2'b11}, // D06.6 (RD = -1)
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0110010111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0110011000, 2'bxx}, // ?
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b00100110, 10'b0110011001, 2'b11}, // D06.1 (RD = -1)
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b10100110, 10'b0110011010, 2'b11}, // D06.5 (RD = -1)
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b00000110, 10'b0110011011, 2'b01}, // D06.0 (RD = -1)
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b01100110, 10'b0110011100, 2'b11}, // D06.3 (RD = -1)
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b10000110, 10'b0110011101, 2'b01}, // D06.4 (RD = -1)
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b11100110, 10'b0110011110, 2'b01}, // D06.7 (RD = -1)
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0110011111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0110100000, 2'bxx}, // ?
    {1'b1, 1'b0, 1'b0, 2'b11, 8'b11110110, 10'b0110100001, 2'b11}, // D22.7 (RD = +1) WRONG RDF
    {1'b1, 1'b0, 1'b0, 2'b11, 8'b10010110, 10'b0110100010, 2'b11}, // D22.4 (RD = +1) WRONG RDF
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0110100011, 2'bxx}, // ?
    {1'b1, 1'b0, 1'b0, 2'b11, 8'b00010110, 10'b0110100100, 2'b11}, // D22.0 (RD = +1) WRONG RDF
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b01010110, 10'b0110100101, 2'b11}, // D22.2 (RD = -1)
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b11010110, 10'b0110100110, 2'b11}, // D22.6 (RD = -1)
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0110100111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0110101000, 2'bxx}, // ?
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b00110110, 10'b0110101001, 2'b11}, // D22.1 (RD = -1)
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b10110110, 10'b0110101010, 2'b11}, // D22.5 (RD = -1)
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b00010110, 10'b0110101011, 2'b01}, // D22.0 (RD = -1)
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b01110110, 10'b0110101100, 2'b11}, // D22.3 (RD = -1)
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b10010110, 10'b0110101101, 2'b01}, // D22.4 (RD = -1)
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b11110110, 10'b0110101110, 2'b01}, // D22.7 (RD = -1)
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0110101111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0110110000, 2'bxx}, // ?
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b11110000, 10'b0110110001, 2'b11}, // D16.7 (RD = -1)
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b10010000, 10'b0110110010, 2'b11}, // D16.4 (RD = -1)
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b01110000, 10'b0110110011, 2'b01}, // D16.3 (RD = -1)
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b00010000, 10'b0110110100, 2'b11}, // D16.0 (RD = -1)
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b01010000, 10'b0110110101, 2'b01}, // D16.2 (RD = -1)
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b11010000, 10'b0110110110, 2'b01}, // D16.6 (RD = -1)
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0110110111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0110111000, 2'bxx}, // ?
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b00110000, 10'b0110111001, 2'b01}, // D16.1 (RD = -1)
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b10110000, 10'b0110111010, 2'b01}, // D16.5 (RD = -1)
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0110111011, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0110111100, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0110111101, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0110111110, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0110111111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0111000000, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0111000001, 2'bxx}, // ?
    {1'b1, 1'b0, 1'b0, 2'b11, 8'b10001110, 10'b0111000010, 2'b11}, // D14.4 (RD = +1) WRONG RDF
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0111000011, 2'bxx}, // ?
    {1'b1, 1'b0, 1'b0, 2'b11, 8'b00001110, 10'b0111000100, 2'b11}, // D14.0 (RD = +1) WRONG RDF
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b01001110, 10'b0111000101, 2'b11}, // D14.2 (RD = -1)
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b11001110, 10'b0111000110, 2'b11}, // D14.6 (RD = -1)
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0111000111, 2'bxx}, // ?
    {1'b1, 1'b0, 1'b0, 2'b11, 8'b11101110, 10'b0111001000, 2'b11}, // D14.7 (RD = +1) WRONG RDF
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b00101110, 10'b0111001001, 2'b11}, // D14.1 (RD = -1)
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b10101110, 10'b0111001010, 2'b11}, // D14.5 (RD = -1)
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b00001110, 10'b0111001011, 2'b01}, // D14.0 (RD = -1)
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b01101110, 10'b0111001100, 2'b11}, // D14.3 (RD = -1)
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b10001110, 10'b0111001101, 2'b01}, // D14.4 (RD = -1)
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b11101110, 10'b0111001110, 2'b01}, // D14.7 (RD = -1)
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0111001111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0111010000, 2'bxx}, // ?
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b11100001, 10'b0111010001, 2'b11}, // D01.7 (RD = -1)
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b10000001, 10'b0111010010, 2'b11}, // D01.4 (RD = -1)
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b01100001, 10'b0111010011, 2'b01}, // D01.3 (RD = -1)
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b00000001, 10'b0111010100, 2'b11}, // D01.0 (RD = -1)
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b01000001, 10'b0111010101, 2'b01}, // D01.2 (RD = -1)
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b11000001, 10'b0111010110, 2'b01}, // D01.6 (RD = -1)
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0111010111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0111011000, 2'bxx}, // ?
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b00100001, 10'b0111011001, 2'b01}, // D01.1 (RD = -1)
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b10100001, 10'b0111011010, 2'b01}, // D01.5 (RD = -1)
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0111011011, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0111011100, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0111011101, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0111011110, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0111011111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0111100000, 2'bxx}, // ?
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b11111110, 10'b0111100001, 2'b11}, // D30.7 (RD = -1)
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b10011110, 10'b0111100010, 2'b11}, // D30.4 (RD = -1)
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b01111110, 10'b0111100011, 2'b01}, // D30.3 (RD = -1)
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b00011110, 10'b0111100100, 2'b11}, // D30.0 (RD = -1)
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b01011110, 10'b0111100101, 2'b01}, // D30.2 (RD = -1)
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b11011110, 10'b0111100110, 2'b01}, // D30.6 (RD = -1)
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0111100111, 2'bxx}, // ?
    {1'b0, 1'b0, 1'b1, 2'b11, 8'b11111110, 10'b0111101000, 2'b11}, // K30.7 (RD = -1)
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b00111110, 10'b0111101001, 2'b01}, // D30.1 (RD = -1)
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b10111110, 10'b0111101010, 2'b01}, // D30.5 (RD = -1)
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0111101011, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0111101100, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0111101101, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0111101110, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0111101111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0111110000, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0111110001, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0111110010, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0111110011, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0111110100, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0111110101, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0111110110, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0111110111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0111111000, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0111111001, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0111111010, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0111111011, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0111111100, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0111111101, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0111111110, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b0111111111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1000000000, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1000000001, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1000000010, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1000000011, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1000000100, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1000000101, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1000000110, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1000000111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1000001000, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1000001001, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1000001010, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1000001011, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1000001100, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1000001101, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1000001110, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1000001111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1000010000, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1000010001, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1000010010, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1000010011, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1000010100, 2'bxx}, // ?
    {1'b1, 1'b0, 1'b0, 2'b11, 8'b01011110, 10'b1000010101, 2'b11}, // D30.2 (RD = +1) WRONG RDF
    {1'b1, 1'b0, 1'b0, 2'b11, 8'b11011110, 10'b1000010110, 2'b11}, // D30.6 (RD = +1) WRONG RDF
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1000010111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1000011000, 2'bxx}, // ?
    {1'b1, 1'b0, 1'b0, 2'b11, 8'b00111110, 10'b1000011001, 2'b11}, // D30.1 (RD = +1) WRONG RDF
    {1'b1, 1'b0, 1'b0, 2'b11, 8'b10111110, 10'b1000011010, 2'b11}, // D30.5 (RD = +1) WRONG RDF
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1000011011, 2'bxx}, // ?
    {1'b1, 1'b0, 1'b0, 2'b11, 8'b01111110, 10'b1000011100, 2'b11}, // D30.3 (RD = +1) WRONG RDF
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1000011101, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1000011110, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1000011111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1000100000, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1000100001, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1000100010, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1000100011, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1000100100, 2'bxx}, // ?
    {1'b1, 1'b0, 1'b0, 2'b11, 8'b01000001, 10'b1000100101, 2'b11}, // D01.2 (RD = +1) WRONG RDF
    {1'b1, 1'b0, 1'b0, 2'b11, 8'b11000001, 10'b1000100110, 2'b11}, // D01.6 (RD = +1) WRONG RDF
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1000100111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1000101000, 2'bxx}, // ?
    {1'b1, 1'b0, 1'b0, 2'b11, 8'b00100001, 10'b1000101001, 2'b11}, // D01.1 (RD = +1) WRONG RDF
    {1'b1, 1'b0, 1'b0, 2'b11, 8'b10100001, 10'b1000101010, 2'b11}, // D01.5 (RD = +1) WRONG RDF
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1000101011, 2'bxx}, // ?
    {1'b1, 1'b0, 1'b0, 2'b11, 8'b01100001, 10'b1000101100, 2'b11}, // D01.3 (RD = +1) WRONG RDF
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1000101101, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1000101110, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1000101111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1000110000, 2'bxx}, // ?
    {1'b1, 1'b0, 1'b0, 2'b11, 8'b11110001, 10'b1000110001, 2'b11}, // D17.7 (RD = +1) WRONG RDF
    {1'b1, 1'b0, 1'b0, 2'b11, 8'b10010001, 10'b1000110010, 2'b11}, // D17.4 (RD = +1) WRONG RDF
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1000110011, 2'bxx}, // ?
    {1'b1, 1'b0, 1'b0, 2'b11, 8'b00010001, 10'b1000110100, 2'b11}, // D17.0 (RD = +1) WRONG RDF
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b01010001, 10'b1000110101, 2'b11}, // D17.2 (RD = -1)
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b11010001, 10'b1000110110, 2'b11}, // D17.6 (RD = -1)
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b11110001, 10'b1000110111, 2'b01}, // D17.7 (RD = -1)
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1000111000, 2'bxx}, // ?
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b00110001, 10'b1000111001, 2'b11}, // D17.1 (RD = -1)
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b10110001, 10'b1000111010, 2'b11}, // D17.5 (RD = -1)
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b00010001, 10'b1000111011, 2'b01}, // D17.0 (RD = -1)
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b01110001, 10'b1000111100, 2'b11}, // D17.3 (RD = -1)
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b10010001, 10'b1000111101, 2'b01}, // D17.4 (RD = -1)
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1000111110, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1000111111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1001000000, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1001000001, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1001000010, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1001000011, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1001000100, 2'bxx}, // ?
    {1'b1, 1'b0, 1'b0, 2'b11, 8'b01010000, 10'b1001000101, 2'b11}, // D16.2 (RD = +1) WRONG RDF
    {1'b1, 1'b0, 1'b0, 2'b11, 8'b11010000, 10'b1001000110, 2'b11}, // D16.6 (RD = +1) WRONG RDF
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1001000111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1001001000, 2'bxx}, // ?
    {1'b1, 1'b0, 1'b0, 2'b11, 8'b00110000, 10'b1001001001, 2'b11}, // D16.1 (RD = +1) WRONG RDF
    {1'b1, 1'b0, 1'b0, 2'b11, 8'b10110000, 10'b1001001010, 2'b11}, // D16.5 (RD = +1) WRONG RDF
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1001001011, 2'bxx}, // ?
    {1'b1, 1'b0, 1'b0, 2'b11, 8'b01110000, 10'b1001001100, 2'b11}, // D16.3 (RD = +1) WRONG RDF
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1001001101, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1001001110, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1001001111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1001010000, 2'bxx}, // ?
    {1'b1, 1'b0, 1'b0, 2'b11, 8'b11101001, 10'b1001010001, 2'b11}, // D09.7 (RD = +1) WRONG RDF
    {1'b1, 1'b0, 1'b0, 2'b11, 8'b10001001, 10'b1001010010, 2'b11}, // D09.4 (RD = +1) WRONG RDF
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1001010011, 2'bxx}, // ?
    {1'b1, 1'b0, 1'b0, 2'b11, 8'b00001001, 10'b1001010100, 2'b11}, // D09.0 (RD = +1) WRONG RDF
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b01001001, 10'b1001010101, 2'b11}, // D09.2 (RD = -1)
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b11001001, 10'b1001010110, 2'b11}, // D09.6 (RD = -1)
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1001010111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1001011000, 2'bxx}, // ?
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b00101001, 10'b1001011001, 2'b11}, // D09.1 (RD = -1)
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b10101001, 10'b1001011010, 2'b11}, // D09.5 (RD = -1)
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b00001001, 10'b1001011011, 2'b01}, // D09.0 (RD = -1)
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b01101001, 10'b1001011100, 2'b11}, // D09.3 (RD = -1)
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b10001001, 10'b1001011101, 2'b01}, // D09.4 (RD = -1)
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b11101001, 10'b1001011110, 2'b01}, // D09.7 (RD = -1)
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1001011111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1001100000, 2'bxx}, // ?
    {1'b1, 1'b0, 1'b0, 2'b11, 8'b11111001, 10'b1001100001, 2'b11}, // D25.7 (RD = +1) WRONG RDF
    {1'b1, 1'b0, 1'b0, 2'b11, 8'b10011001, 10'b1001100010, 2'b11}, // D25.4 (RD = +1) WRONG RDF
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1001100011, 2'bxx}, // ?
    {1'b1, 1'b0, 1'b0, 2'b11, 8'b00011001, 10'b1001100100, 2'b11}, // D25.0 (RD = +1) WRONG RDF
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b01011001, 10'b1001100101, 2'b11}, // D25.2 (RD = -1)
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b11011001, 10'b1001100110, 2'b11}, // D25.6 (RD = -1)
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1001100111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1001101000, 2'bxx}, // ?
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b00111001, 10'b1001101001, 2'b11}, // D25.1 (RD = -1)
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b10111001, 10'b1001101010, 2'b11}, // D25.5 (RD = -1)
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b00011001, 10'b1001101011, 2'b01}, // D25.0 (RD = -1)
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b01111001, 10'b1001101100, 2'b11}, // D25.3 (RD = -1)
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b10011001, 10'b1001101101, 2'b01}, // D25.4 (RD = -1)
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b11111001, 10'b1001101110, 2'b01}, // D25.7 (RD = -1)
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1001101111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1001110000, 2'bxx}, // ?
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b11100000, 10'b1001110001, 2'b11}, // D00.7 (RD = -1)
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b10000000, 10'b1001110010, 2'b11}, // D00.4 (RD = -1)
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b01100000, 10'b1001110011, 2'b01}, // D00.3 (RD = -1)
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b00000000, 10'b1001110100, 2'b11}, // D00.0 (RD = -1)
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b01000000, 10'b1001110101, 2'b01}, // D00.2 (RD = -1)
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b11000000, 10'b1001110110, 2'b01}, // D00.6 (RD = -1)
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1001110111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1001111000, 2'bxx}, // ?
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b00100000, 10'b1001111001, 2'b01}, // D00.1 (RD = -1)
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b10100000, 10'b1001111010, 2'b01}, // D00.5 (RD = -1)
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1001111011, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1001111100, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1001111101, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1001111110, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1001111111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1010000000, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1010000001, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1010000010, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1010000011, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1010000100, 2'bxx}, // ?
    {1'b1, 1'b0, 1'b0, 2'b11, 8'b01001111, 10'b1010000101, 2'b11}, // D15.2 (RD = +1) WRONG RDF
    {1'b1, 1'b0, 1'b0, 2'b11, 8'b11001111, 10'b1010000110, 2'b11}, // D15.6 (RD = +1) WRONG RDF
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1010000111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1010001000, 2'bxx}, // ?
    {1'b1, 1'b0, 1'b0, 2'b11, 8'b00101111, 10'b1010001001, 2'b11}, // D15.1 (RD = +1) WRONG RDF
    {1'b1, 1'b0, 1'b0, 2'b11, 8'b10101111, 10'b1010001010, 2'b11}, // D15.5 (RD = +1) WRONG RDF
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1010001011, 2'bxx}, // ?
    {1'b1, 1'b0, 1'b0, 2'b11, 8'b01101111, 10'b1010001100, 2'b11}, // D15.3 (RD = +1) WRONG RDF
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1010001101, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1010001110, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1010001111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1010010000, 2'bxx}, // ?
    {1'b1, 1'b0, 1'b0, 2'b11, 8'b11100101, 10'b1010010001, 2'b11}, // D05.7 (RD = +1) WRONG RDF
    {1'b1, 1'b0, 1'b0, 2'b11, 8'b10000101, 10'b1010010010, 2'b11}, // D05.4 (RD = +1) WRONG RDF
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1010010011, 2'bxx}, // ?
    {1'b1, 1'b0, 1'b0, 2'b11, 8'b00000101, 10'b1010010100, 2'b11}, // D05.0 (RD = +1) WRONG RDF
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b01000101, 10'b1010010101, 2'b11}, // D05.2 (RD = -1)
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b11000101, 10'b1010010110, 2'b11}, // D05.6 (RD = -1)
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1010010111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1010011000, 2'bxx}, // ?
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b00100101, 10'b1010011001, 2'b11}, // D05.1 (RD = -1)
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b10100101, 10'b1010011010, 2'b11}, // D05.5 (RD = -1)
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b00000101, 10'b1010011011, 2'b01}, // D05.0 (RD = -1)
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b01100101, 10'b1010011100, 2'b11}, // D05.3 (RD = -1)
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b10000101, 10'b1010011101, 2'b01}, // D05.4 (RD = -1)
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b11100101, 10'b1010011110, 2'b01}, // D05.7 (RD = -1)
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1010011111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1010100000, 2'bxx}, // ?
    {1'b1, 1'b0, 1'b0, 2'b11, 8'b11110101, 10'b1010100001, 2'b11}, // D21.7 (RD = +1) WRONG RDF
    {1'b1, 1'b0, 1'b0, 2'b11, 8'b10010101, 10'b1010100010, 2'b11}, // D21.4 (RD = +1) WRONG RDF
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1010100011, 2'bxx}, // ?
    {1'b1, 1'b0, 1'b0, 2'b11, 8'b00010101, 10'b1010100100, 2'b11}, // D21.0 (RD = +1) WRONG RDF
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b01010101, 10'b1010100101, 2'b11}, // D21.2 (RD = -1)
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b11010101, 10'b1010100110, 2'b11}, // D21.6 (RD = -1)
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1010100111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1010101000, 2'bxx}, // ?
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b00110101, 10'b1010101001, 2'b11}, // D21.1 (RD = -1)
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b10110101, 10'b1010101010, 2'b11}, // D21.5 (RD = -1)
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b00010101, 10'b1010101011, 2'b01}, // D21.0 (RD = -1)
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b01110101, 10'b1010101100, 2'b11}, // D21.3 (RD = -1)
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b10010101, 10'b1010101101, 2'b01}, // D21.4 (RD = -1)
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b11110101, 10'b1010101110, 2'b01}, // D21.7 (RD = -1)
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1010101111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1010110000, 2'bxx}, // ?
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b11111111, 10'b1010110001, 2'b11}, // D31.7 (RD = -1)
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b10011111, 10'b1010110010, 2'b11}, // D31.4 (RD = -1)
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b01111111, 10'b1010110011, 2'b01}, // D31.3 (RD = -1)
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b00011111, 10'b1010110100, 2'b11}, // D31.0 (RD = -1)
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b01011111, 10'b1010110101, 2'b01}, // D31.2 (RD = -1)
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b11011111, 10'b1010110110, 2'b01}, // D31.6 (RD = -1)
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1010110111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1010111000, 2'bxx}, // ?
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b00111111, 10'b1010111001, 2'b01}, // D31.1 (RD = -1)
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b10111111, 10'b1010111010, 2'b01}, // D31.5 (RD = -1)
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1010111011, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1010111100, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1010111101, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1010111110, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1010111111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1011000000, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1011000001, 2'bxx}, // ?
    {1'b1, 1'b0, 1'b0, 2'b11, 8'b10001101, 10'b1011000010, 2'b11}, // D13.4 (RD = +1) WRONG RDF
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1011000011, 2'bxx}, // ?
    {1'b1, 1'b0, 1'b0, 2'b11, 8'b00001101, 10'b1011000100, 2'b11}, // D13.0 (RD = +1) WRONG RDF
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b01001101, 10'b1011000101, 2'b11}, // D13.2 (RD = -1)
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b11001101, 10'b1011000110, 2'b11}, // D13.6 (RD = -1)
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1011000111, 2'bxx}, // ?
    {1'b1, 1'b0, 1'b0, 2'b11, 8'b11101101, 10'b1011001000, 2'b11}, // D13.7 (RD = +1) WRONG RDF
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b00101101, 10'b1011001001, 2'b11}, // D13.1 (RD = -1)
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b10101101, 10'b1011001010, 2'b11}, // D13.5 (RD = -1)
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b00001101, 10'b1011001011, 2'b01}, // D13.0 (RD = -1)
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b01101101, 10'b1011001100, 2'b11}, // D13.3 (RD = -1)
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b10001101, 10'b1011001101, 2'b01}, // D13.4 (RD = -1)
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b11101101, 10'b1011001110, 2'b01}, // D13.7 (RD = -1)
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1011001111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1011010000, 2'bxx}, // ?
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b11100010, 10'b1011010001, 2'b11}, // D02.7 (RD = -1)
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b10000010, 10'b1011010010, 2'b11}, // D02.4 (RD = -1)
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b01100010, 10'b1011010011, 2'b01}, // D02.3 (RD = -1)
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b00000010, 10'b1011010100, 2'b11}, // D02.0 (RD = -1)
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b01000010, 10'b1011010101, 2'b01}, // D02.2 (RD = -1)
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b11000010, 10'b1011010110, 2'b01}, // D02.6 (RD = -1)
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1011010111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1011011000, 2'bxx}, // ?
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b00100010, 10'b1011011001, 2'b01}, // D02.1 (RD = -1)
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b10100010, 10'b1011011010, 2'b01}, // D02.5 (RD = -1)
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1011011011, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1011011100, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1011011101, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1011011110, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1011011111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1011100000, 2'bxx}, // ?
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b11111101, 10'b1011100001, 2'b11}, // D29.7 (RD = -1)
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b10011101, 10'b1011100010, 2'b11}, // D29.4 (RD = -1)
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b01111101, 10'b1011100011, 2'b01}, // D29.3 (RD = -1)
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b00011101, 10'b1011100100, 2'b11}, // D29.0 (RD = -1)
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b01011101, 10'b1011100101, 2'b01}, // D29.2 (RD = -1)
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b11011101, 10'b1011100110, 2'b01}, // D29.6 (RD = -1)
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1011100111, 2'bxx}, // ?
    {1'b0, 1'b0, 1'b1, 2'b11, 8'b11111101, 10'b1011101000, 2'b11}, // K29.7 (RD = -1)
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b00111101, 10'b1011101001, 2'b01}, // D29.1 (RD = -1)
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b10111101, 10'b1011101010, 2'b01}, // D29.5 (RD = -1)
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1011101011, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1011101100, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1011101101, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1011101110, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1011101111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1011110000, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1011110001, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1011110010, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1011110011, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1011110100, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1011110101, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1011110110, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1011110111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1011111000, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1011111001, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1011111010, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1011111011, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1011111100, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1011111101, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1011111110, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1011111111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1100000000, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1100000001, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1100000010, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1100000011, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1100000100, 2'bxx}, // ?
    {1'b1, 1'b0, 1'b1, 2'b11, 8'b10111100, 10'b1100000101, 2'b11}, // K28.5 (RD = +1) WRONG RDF
    {1'b1, 1'b0, 1'b1, 2'b11, 8'b00111100, 10'b1100000110, 2'b11}, // K28.1 (RD = +1) WRONG RDF
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1100000111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1100001000, 2'bxx}, // ?
    {1'b1, 1'b0, 1'b1, 2'b11, 8'b11011100, 10'b1100001001, 2'b11}, // K28.6 (RD = +1) WRONG RDF
    {1'b1, 1'b0, 1'b1, 2'b11, 8'b01011100, 10'b1100001010, 2'b11}, // K28.2 (RD = +1) WRONG RDF
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1100001011, 2'bxx}, // ?
    {1'b1, 1'b0, 1'b1, 2'b11, 8'b01111100, 10'b1100001100, 2'b11}, // K28.3 (RD = +1) WRONG RDF
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1100001101, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1100001110, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1100001111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1100010000, 2'bxx}, // ?
    {1'b1, 1'b0, 1'b0, 2'b11, 8'b11100011, 10'b1100010001, 2'b11}, // D03.7 (RD = +1) WRONG RDF
    {1'b1, 1'b0, 1'b0, 2'b11, 8'b10000011, 10'b1100010010, 2'b11}, // D03.4 (RD = +1) WRONG RDF
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1100010011, 2'bxx}, // ?
    {1'b1, 1'b0, 1'b0, 2'b11, 8'b00000011, 10'b1100010100, 2'b11}, // D03.0 (RD = +1) WRONG RDF
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b01000011, 10'b1100010101, 2'b11}, // D03.2 (RD = -1)
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b11000011, 10'b1100010110, 2'b11}, // D03.6 (RD = -1)
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1100010111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1100011000, 2'bxx}, // ?
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b00100011, 10'b1100011001, 2'b11}, // D03.1 (RD = -1)
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b10100011, 10'b1100011010, 2'b11}, // D03.5 (RD = -1)
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b00000011, 10'b1100011011, 2'b01}, // D03.0 (RD = -1)
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b01100011, 10'b1100011100, 2'b11}, // D03.3 (RD = -1)
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b10000011, 10'b1100011101, 2'b01}, // D03.4 (RD = -1)
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b11100011, 10'b1100011110, 2'b01}, // D03.7 (RD = -1)
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1100011111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1100100000, 2'bxx}, // ?
    {1'b1, 1'b0, 1'b0, 2'b11, 8'b11110011, 10'b1100100001, 2'b11}, // D19.7 (RD = +1) WRONG RDF
    {1'b1, 1'b0, 1'b0, 2'b11, 8'b10010011, 10'b1100100010, 2'b11}, // D19.4 (RD = +1) WRONG RDF
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1100100011, 2'bxx}, // ?
    {1'b1, 1'b0, 1'b0, 2'b11, 8'b00010011, 10'b1100100100, 2'b11}, // D19.0 (RD = +1) WRONG RDF
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b01010011, 10'b1100100101, 2'b11}, // D19.2 (RD = -1)
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b11010011, 10'b1100100110, 2'b11}, // D19.6 (RD = -1)
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1100100111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1100101000, 2'bxx}, // ?
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b00110011, 10'b1100101001, 2'b11}, // D19.1 (RD = -1)
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b10110011, 10'b1100101010, 2'b11}, // D19.5 (RD = -1)
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b00010011, 10'b1100101011, 2'b01}, // D19.0 (RD = -1)
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b01110011, 10'b1100101100, 2'b11}, // D19.3 (RD = -1)
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b10010011, 10'b1100101101, 2'b01}, // D19.4 (RD = -1)
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b11110011, 10'b1100101110, 2'b01}, // D19.7 (RD = -1)
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1100101111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1100110000, 2'bxx}, // ?
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b11111000, 10'b1100110001, 2'b11}, // D24.7 (RD = -1)
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b10011000, 10'b1100110010, 2'b11}, // D24.4 (RD = -1)
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b01111000, 10'b1100110011, 2'b01}, // D24.3 (RD = -1)
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b00011000, 10'b1100110100, 2'b11}, // D24.0 (RD = -1)
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b01011000, 10'b1100110101, 2'b01}, // D24.2 (RD = -1)
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b11011000, 10'b1100110110, 2'b01}, // D24.6 (RD = -1)
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1100110111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1100111000, 2'bxx}, // ?
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b00111000, 10'b1100111001, 2'b01}, // D24.1 (RD = -1)
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b10111000, 10'b1100111010, 2'b01}, // D24.5 (RD = -1)
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1100111011, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1100111100, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1100111101, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1100111110, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1100111111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1101000000, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1101000001, 2'bxx}, // ?
    {1'b1, 1'b0, 1'b0, 2'b11, 8'b10001011, 10'b1101000010, 2'b11}, // D11.4 (RD = +1) WRONG RDF
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1101000011, 2'bxx}, // ?
    {1'b1, 1'b0, 1'b0, 2'b11, 8'b00001011, 10'b1101000100, 2'b11}, // D11.0 (RD = +1) WRONG RDF
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b01001011, 10'b1101000101, 2'b11}, // D11.2 (RD = -1)
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b11001011, 10'b1101000110, 2'b11}, // D11.6 (RD = -1)
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1101000111, 2'bxx}, // ?
    {1'b1, 1'b0, 1'b0, 2'b11, 8'b11101011, 10'b1101001000, 2'b11}, // D11.7 (RD = +1) WRONG RDF
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b00101011, 10'b1101001001, 2'b11}, // D11.1 (RD = -1)
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b10101011, 10'b1101001010, 2'b11}, // D11.5 (RD = -1)
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b00001011, 10'b1101001011, 2'b01}, // D11.0 (RD = -1)
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b01101011, 10'b1101001100, 2'b11}, // D11.3 (RD = -1)
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b10001011, 10'b1101001101, 2'b01}, // D11.4 (RD = -1)
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b11101011, 10'b1101001110, 2'b01}, // D11.7 (RD = -1)
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1101001111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1101010000, 2'bxx}, // ?
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b11100100, 10'b1101010001, 2'b11}, // D04.7 (RD = -1)
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b10000100, 10'b1101010010, 2'b11}, // D04.4 (RD = -1)
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b01100100, 10'b1101010011, 2'b01}, // D04.3 (RD = -1)
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b00000100, 10'b1101010100, 2'b11}, // D04.0 (RD = -1)
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b01000100, 10'b1101010101, 2'b01}, // D04.2 (RD = -1)
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b11000100, 10'b1101010110, 2'b01}, // D04.6 (RD = -1)
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1101010111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1101011000, 2'bxx}, // ?
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b00100100, 10'b1101011001, 2'b01}, // D04.1 (RD = -1)
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b10100100, 10'b1101011010, 2'b01}, // D04.5 (RD = -1)
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1101011011, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1101011100, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1101011101, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1101011110, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1101011111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1101100000, 2'bxx}, // ?
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b11111011, 10'b1101100001, 2'b11}, // D27.7 (RD = -1)
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b10011011, 10'b1101100010, 2'b11}, // D27.4 (RD = -1)
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b01111011, 10'b1101100011, 2'b01}, // D27.3 (RD = -1)
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b00011011, 10'b1101100100, 2'b11}, // D27.0 (RD = -1)
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b01011011, 10'b1101100101, 2'b01}, // D27.2 (RD = -1)
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b11011011, 10'b1101100110, 2'b01}, // D27.6 (RD = -1)
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1101100111, 2'bxx}, // ?
    {1'b0, 1'b0, 1'b1, 2'b11, 8'b11111011, 10'b1101101000, 2'b11}, // K27.7 (RD = -1)
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b00111011, 10'b1101101001, 2'b01}, // D27.1 (RD = -1)
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b10111011, 10'b1101101010, 2'b01}, // D27.5 (RD = -1)
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1101101011, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1101101100, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1101101101, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1101101110, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1101101111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1101110000, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1101110001, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1101110010, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1101110011, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1101110100, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1101110101, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1101110110, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1101110111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1101111000, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1101111001, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1101111010, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1101111011, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1101111100, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1101111101, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1101111110, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1101111111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1110000000, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1110000001, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1110000010, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1110000011, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1110000100, 2'bxx}, // ?
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b01000111, 10'b1110000101, 2'b11}, // D07.2 (RD = -1)
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b11000111, 10'b1110000110, 2'b11}, // D07.6 (RD = -1)
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1110000111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1110001000, 2'bxx}, // ?
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b00100111, 10'b1110001001, 2'b11}, // D07.1 (RD = -1)
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b10100111, 10'b1110001010, 2'b11}, // D07.5 (RD = -1)
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b00000111, 10'b1110001011, 2'b01}, // D07.0 (RD = -1)
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b01100111, 10'b1110001100, 2'b11}, // D07.3 (RD = -1)
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b10000111, 10'b1110001101, 2'b01}, // D07.4 (RD = -1)
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b11100111, 10'b1110001110, 2'b01}, // D07.7 (RD = -1)
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1110001111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1110010000, 2'bxx}, // ?
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b11101000, 10'b1110010001, 2'b11}, // D08.7 (RD = -1)
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b10001000, 10'b1110010010, 2'b11}, // D08.4 (RD = -1)
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b01101000, 10'b1110010011, 2'b01}, // D08.3 (RD = -1)
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b00001000, 10'b1110010100, 2'b11}, // D08.0 (RD = -1)
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b01001000, 10'b1110010101, 2'b01}, // D08.2 (RD = -1)
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b11001000, 10'b1110010110, 2'b01}, // D08.6 (RD = -1)
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1110010111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1110011000, 2'bxx}, // ?
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b00101000, 10'b1110011001, 2'b01}, // D08.1 (RD = -1)
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b10101000, 10'b1110011010, 2'b01}, // D08.5 (RD = -1)
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1110011011, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1110011100, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1110011101, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1110011110, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1110011111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1110100000, 2'bxx}, // ?
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b11110111, 10'b1110100001, 2'b11}, // D23.7 (RD = -1)
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b10010111, 10'b1110100010, 2'b11}, // D23.4 (RD = -1)
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b01110111, 10'b1110100011, 2'b01}, // D23.3 (RD = -1)
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b00010111, 10'b1110100100, 2'b11}, // D23.0 (RD = -1)
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b01010111, 10'b1110100101, 2'b01}, // D23.2 (RD = -1)
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b11010111, 10'b1110100110, 2'b01}, // D23.6 (RD = -1)
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1110100111, 2'bxx}, // ?
    {1'b0, 1'b0, 1'b1, 2'b11, 8'b11110111, 10'b1110101000, 2'b11}, // K23.7 (RD = -1)
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b00110111, 10'b1110101001, 2'b01}, // D23.1 (RD = -1)
    {1'b0, 1'b0, 1'b0, 2'b11, 8'b10110111, 10'b1110101010, 2'b01}, // D23.5 (RD = -1)
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1110101011, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1110101100, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1110101101, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1110101110, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1110101111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1110110000, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1110110001, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1110110010, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1110110011, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1110110100, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1110110101, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1110110110, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1110110111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1110111000, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1110111001, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1110111010, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1110111011, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1110111100, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1110111101, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1110111110, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1110111111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1111000000, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1111000001, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1111000010, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1111000011, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1111000100, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1111000101, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1111000110, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1111000111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1111001000, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1111001001, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1111001010, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1111001011, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1111001100, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1111001101, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1111001110, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1111001111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1111010000, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1111010001, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1111010010, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1111010011, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1111010100, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1111010101, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1111010110, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1111010111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1111011000, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1111011001, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1111011010, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1111011011, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1111011100, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1111011101, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1111011110, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1111011111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1111100000, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1111100001, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1111100010, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1111100011, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1111100100, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1111100101, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1111100110, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1111100111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1111101000, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1111101001, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1111101010, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1111101011, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1111101100, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1111101101, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1111101110, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1111101111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1111110000, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1111110001, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1111110010, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1111110011, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1111110100, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1111110101, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1111110110, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1111110111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1111111000, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1111111001, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1111111010, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1111111011, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1111111100, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1111111101, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1111111110, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b11, 8'bxxxxxxxx, 10'b1111111111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0000000000, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0000000001, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0000000010, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0000000011, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0000000100, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0000000101, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0000000110, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0000000111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0000001000, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0000001001, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0000001010, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0000001011, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0000001100, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0000001101, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0000001110, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0000001111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0000010000, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0000010001, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0000010010, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0000010011, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0000010100, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0000010101, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0000010110, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0000010111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0000011000, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0000011001, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0000011010, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0000011011, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0000011100, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0000011101, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0000011110, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0000011111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0000100000, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0000100001, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0000100010, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0000100011, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0000100100, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0000100101, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0000100110, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0000100111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0000101000, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0000101001, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0000101010, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0000101011, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0000101100, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0000101101, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0000101110, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0000101111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0000110000, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0000110001, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0000110010, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0000110011, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0000110100, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0000110101, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0000110110, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0000110111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0000111000, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0000111001, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0000111010, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0000111011, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0000111100, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0000111101, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0000111110, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0000111111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0001000000, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0001000001, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0001000010, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0001000011, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0001000100, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0001000101, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0001000110, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0001000111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0001001000, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0001001001, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0001001010, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0001001011, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0001001100, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0001001101, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0001001110, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0001001111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0001010000, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0001010001, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0001010010, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0001010011, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0001010100, 2'bxx}, // ?
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b01010111, 10'b0001010101, 2'b11}, // D23.2 (RD = +1)
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b11010111, 10'b0001010110, 2'b11}, // D23.6 (RD = +1)
    {1'b0, 1'b0, 1'b1, 2'b01, 8'b11110111, 10'b0001010111, 2'b01}, // K23.7 (RD = +1)
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0001011000, 2'bxx}, // ?
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b00110111, 10'b0001011001, 2'b11}, // D23.1 (RD = +1)
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b10110111, 10'b0001011010, 2'b11}, // D23.5 (RD = +1)
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b00010111, 10'b0001011011, 2'b01}, // D23.0 (RD = +1)
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b01110111, 10'b0001011100, 2'b11}, // D23.3 (RD = +1)
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b10010111, 10'b0001011101, 2'b01}, // D23.4 (RD = +1)
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b11110111, 10'b0001011110, 2'b01}, // D23.7 (RD = +1)
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0001011111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0001100000, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0001100001, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0001100010, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0001100011, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0001100100, 2'bxx}, // ?
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b01001000, 10'b0001100101, 2'b11}, // D08.2 (RD = +1)
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b11001000, 10'b0001100110, 2'b11}, // D08.6 (RD = +1)
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0001100111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0001101000, 2'bxx}, // ?
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b00101000, 10'b0001101001, 2'b11}, // D08.1 (RD = +1)
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b10101000, 10'b0001101010, 2'b11}, // D08.5 (RD = +1)
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b00001000, 10'b0001101011, 2'b01}, // D08.0 (RD = +1)
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b01101000, 10'b0001101100, 2'b11}, // D08.3 (RD = +1)
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b10001000, 10'b0001101101, 2'b01}, // D08.4 (RD = +1)
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b11101000, 10'b0001101110, 2'b01}, // D08.7 (RD = +1)
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0001101111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0001110000, 2'bxx}, // ?
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b11100111, 10'b0001110001, 2'b11}, // D07.7 (RD = +1)
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b10000111, 10'b0001110010, 2'b11}, // D07.4 (RD = +1)
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b01100111, 10'b0001110011, 2'b01}, // D07.3 (RD = +1)
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b00000111, 10'b0001110100, 2'b11}, // D07.0 (RD = +1)
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b01000111, 10'b0001110101, 2'b01}, // D07.2 (RD = +1)
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b11000111, 10'b0001110110, 2'b01}, // D07.6 (RD = +1)
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0001110111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0001111000, 2'bxx}, // ?
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b00100111, 10'b0001111001, 2'b01}, // D07.1 (RD = +1)
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b10100111, 10'b0001111010, 2'b01}, // D07.5 (RD = +1)
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0001111011, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0001111100, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0001111101, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0001111110, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0001111111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0010000000, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0010000001, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0010000010, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0010000011, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0010000100, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0010000101, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0010000110, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0010000111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0010001000, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0010001001, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0010001010, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0010001011, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0010001100, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0010001101, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0010001110, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0010001111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0010010000, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0010010001, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0010010010, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0010010011, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0010010100, 2'bxx}, // ?
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b01011011, 10'b0010010101, 2'b11}, // D27.2 (RD = +1)
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b11011011, 10'b0010010110, 2'b11}, // D27.6 (RD = +1)
    {1'b0, 1'b0, 1'b1, 2'b01, 8'b11111011, 10'b0010010111, 2'b01}, // K27.7 (RD = +1)
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0010011000, 2'bxx}, // ?
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b00111011, 10'b0010011001, 2'b11}, // D27.1 (RD = +1)
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b10111011, 10'b0010011010, 2'b11}, // D27.5 (RD = +1)
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b00011011, 10'b0010011011, 2'b01}, // D27.0 (RD = +1)
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b01111011, 10'b0010011100, 2'b11}, // D27.3 (RD = +1)
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b10011011, 10'b0010011101, 2'b01}, // D27.4 (RD = +1)
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b11111011, 10'b0010011110, 2'b01}, // D27.7 (RD = +1)
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0010011111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0010100000, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0010100001, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0010100010, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0010100011, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0010100100, 2'bxx}, // ?
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b01000100, 10'b0010100101, 2'b11}, // D04.2 (RD = +1)
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b11000100, 10'b0010100110, 2'b11}, // D04.6 (RD = +1)
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0010100111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0010101000, 2'bxx}, // ?
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b00100100, 10'b0010101001, 2'b11}, // D04.1 (RD = +1)
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b10100100, 10'b0010101010, 2'b11}, // D04.5 (RD = +1)
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b00000100, 10'b0010101011, 2'b01}, // D04.0 (RD = +1)
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b01100100, 10'b0010101100, 2'b11}, // D04.3 (RD = +1)
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b10000100, 10'b0010101101, 2'b01}, // D04.4 (RD = +1)
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b11100100, 10'b0010101110, 2'b01}, // D04.7 (RD = +1)
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0010101111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0010110000, 2'bxx}, // ?
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b11110100, 10'b0010110001, 2'b11}, // D20.7 (RD = +1)
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b10010100, 10'b0010110010, 2'b11}, // D20.4 (RD = +1)
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b01110100, 10'b0010110011, 2'b01}, // D20.3 (RD = +1)
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b00010100, 10'b0010110100, 2'b11}, // D20.0 (RD = +1)
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b01010100, 10'b0010110101, 2'b01}, // D20.2 (RD = +1)
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b11010100, 10'b0010110110, 2'b01}, // D20.6 (RD = +1)
    {1'b1, 1'b0, 1'b0, 2'b01, 8'b11110100, 10'b0010110111, 2'b01}, // D20.7 (RD = -1) WRONG RDF
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0010111000, 2'bxx}, // ?
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b00110100, 10'b0010111001, 2'b01}, // D20.1 (RD = +1)
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b10110100, 10'b0010111010, 2'b01}, // D20.5 (RD = +1)
    {1'b1, 1'b0, 1'b0, 2'b01, 8'b00010100, 10'b0010111011, 2'b01}, // D20.0 (RD = -1) WRONG RDF
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0010111100, 2'bxx}, // ?
    {1'b1, 1'b0, 1'b0, 2'b01, 8'b10010100, 10'b0010111101, 2'b01}, // D20.4 (RD = -1) WRONG RDF
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0010111110, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0010111111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0011000000, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0011000001, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0011000010, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0011000011, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0011000100, 2'bxx}, // ?
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b01011000, 10'b0011000101, 2'b11}, // D24.2 (RD = +1)
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b11011000, 10'b0011000110, 2'b11}, // D24.6 (RD = +1)
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0011000111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0011001000, 2'bxx}, // ?
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b00111000, 10'b0011001001, 2'b11}, // D24.1 (RD = +1)
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b10111000, 10'b0011001010, 2'b11}, // D24.5 (RD = +1)
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b00011000, 10'b0011001011, 2'b01}, // D24.0 (RD = +1)
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b01111000, 10'b0011001100, 2'b11}, // D24.3 (RD = +1)
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b10011000, 10'b0011001101, 2'b01}, // D24.4 (RD = +1)
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b11111000, 10'b0011001110, 2'b01}, // D24.7 (RD = +1)
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0011001111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0011010000, 2'bxx}, // ?
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b11101100, 10'b0011010001, 2'b11}, // D12.7 (RD = +1)
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b10001100, 10'b0011010010, 2'b11}, // D12.4 (RD = +1)
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b01101100, 10'b0011010011, 2'b01}, // D12.3 (RD = +1)
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b00001100, 10'b0011010100, 2'b11}, // D12.0 (RD = +1)
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b01001100, 10'b0011010101, 2'b01}, // D12.2 (RD = +1)
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b11001100, 10'b0011010110, 2'b01}, // D12.6 (RD = +1)
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0011010111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0011011000, 2'bxx}, // ?
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b00101100, 10'b0011011001, 2'b01}, // D12.1 (RD = +1)
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b10101100, 10'b0011011010, 2'b01}, // D12.5 (RD = +1)
    {1'b1, 1'b0, 1'b0, 2'b01, 8'b00001100, 10'b0011011011, 2'b01}, // D12.0 (RD = -1) WRONG RDF
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0011011100, 2'bxx}, // ?
    {1'b1, 1'b0, 1'b0, 2'b01, 8'b10001100, 10'b0011011101, 2'b01}, // D12.4 (RD = -1) WRONG RDF
    {1'b1, 1'b0, 1'b0, 2'b01, 8'b11101100, 10'b0011011110, 2'b01}, // D12.7 (RD = -1) WRONG RDF
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0011011111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0011100000, 2'bxx}, // ?
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b11111100, 10'b0011100001, 2'b11}, // D28.7 (RD = +1)
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b10011100, 10'b0011100010, 2'b11}, // D28.4 (RD = +1)
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b01111100, 10'b0011100011, 2'b01}, // D28.3 (RD = +1)
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b00011100, 10'b0011100100, 2'b11}, // D28.0 (RD = +1)
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b01011100, 10'b0011100101, 2'b01}, // D28.2 (RD = +1)
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b11011100, 10'b0011100110, 2'b01}, // D28.6 (RD = +1)
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0011100111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0011101000, 2'bxx}, // ?
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b00111100, 10'b0011101001, 2'b01}, // D28.1 (RD = +1)
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b10111100, 10'b0011101010, 2'b01}, // D28.5 (RD = +1)
    {1'b1, 1'b0, 1'b0, 2'b01, 8'b00011100, 10'b0011101011, 2'b01}, // D28.0 (RD = -1) WRONG RDF
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0011101100, 2'bxx}, // ?
    {1'b1, 1'b0, 1'b0, 2'b01, 8'b10011100, 10'b0011101101, 2'b01}, // D28.4 (RD = -1) WRONG RDF
    {1'b1, 1'b0, 1'b0, 2'b01, 8'b11111100, 10'b0011101110, 2'b01}, // D28.7 (RD = -1) WRONG RDF
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0011101111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0011110000, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0011110001, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0011110010, 2'bxx}, // ?
    {1'b1, 1'b0, 1'b1, 2'b01, 8'b01111100, 10'b0011110011, 2'b01}, // K28.3 (RD = -1) WRONG RDF
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0011110100, 2'bxx}, // ?
    {1'b1, 1'b0, 1'b1, 2'b01, 8'b01011100, 10'b0011110101, 2'b01}, // K28.2 (RD = -1) WRONG RDF
    {1'b1, 1'b0, 1'b1, 2'b01, 8'b11011100, 10'b0011110110, 2'b01}, // K28.6 (RD = -1) WRONG RDF
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0011110111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0011111000, 2'bxx}, // ?
    {1'b1, 1'b0, 1'b1, 2'b01, 8'b00111100, 10'b0011111001, 2'b01}, // K28.1 (RD = -1) WRONG RDF
    {1'b1, 1'b0, 1'b1, 2'b01, 8'b10111100, 10'b0011111010, 2'b01}, // K28.5 (RD = -1) WRONG RDF
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0011111011, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0011111100, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0011111101, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0011111110, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0011111111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0100000000, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0100000001, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0100000010, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0100000011, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0100000100, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0100000101, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0100000110, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0100000111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0100001000, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0100001001, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0100001010, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0100001011, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0100001100, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0100001101, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0100001110, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0100001111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0100010000, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0100010001, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0100010010, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0100010011, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0100010100, 2'bxx}, // ?
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b01011101, 10'b0100010101, 2'b11}, // D29.2 (RD = +1)
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b11011101, 10'b0100010110, 2'b11}, // D29.6 (RD = +1)
    {1'b0, 1'b0, 1'b1, 2'b01, 8'b11111101, 10'b0100010111, 2'b01}, // K29.7 (RD = +1)
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0100011000, 2'bxx}, // ?
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b00111101, 10'b0100011001, 2'b11}, // D29.1 (RD = +1)
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b10111101, 10'b0100011010, 2'b11}, // D29.5 (RD = +1)
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b00011101, 10'b0100011011, 2'b01}, // D29.0 (RD = +1)
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b01111101, 10'b0100011100, 2'b11}, // D29.3 (RD = +1)
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b10011101, 10'b0100011101, 2'b01}, // D29.4 (RD = +1)
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b11111101, 10'b0100011110, 2'b01}, // D29.7 (RD = +1)
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0100011111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0100100000, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0100100001, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0100100010, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0100100011, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0100100100, 2'bxx}, // ?
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b01000010, 10'b0100100101, 2'b11}, // D02.2 (RD = +1)
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b11000010, 10'b0100100110, 2'b11}, // D02.6 (RD = +1)
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0100100111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0100101000, 2'bxx}, // ?
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b00100010, 10'b0100101001, 2'b11}, // D02.1 (RD = +1)
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b10100010, 10'b0100101010, 2'b11}, // D02.5 (RD = +1)
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b00000010, 10'b0100101011, 2'b01}, // D02.0 (RD = +1)
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b01100010, 10'b0100101100, 2'b11}, // D02.3 (RD = +1)
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b10000010, 10'b0100101101, 2'b01}, // D02.4 (RD = +1)
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b11100010, 10'b0100101110, 2'b01}, // D02.7 (RD = +1)
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0100101111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0100110000, 2'bxx}, // ?
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b11110010, 10'b0100110001, 2'b11}, // D18.7 (RD = +1)
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b10010010, 10'b0100110010, 2'b11}, // D18.4 (RD = +1)
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b01110010, 10'b0100110011, 2'b01}, // D18.3 (RD = +1)
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b00010010, 10'b0100110100, 2'b11}, // D18.0 (RD = +1)
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b01010010, 10'b0100110101, 2'b01}, // D18.2 (RD = +1)
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b11010010, 10'b0100110110, 2'b01}, // D18.6 (RD = +1)
    {1'b1, 1'b0, 1'b0, 2'b01, 8'b11110010, 10'b0100110111, 2'b01}, // D18.7 (RD = -1) WRONG RDF
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0100111000, 2'bxx}, // ?
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b00110010, 10'b0100111001, 2'b01}, // D18.1 (RD = +1)
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b10110010, 10'b0100111010, 2'b01}, // D18.5 (RD = +1)
    {1'b1, 1'b0, 1'b0, 2'b01, 8'b00010010, 10'b0100111011, 2'b01}, // D18.0 (RD = -1) WRONG RDF
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0100111100, 2'bxx}, // ?
    {1'b1, 1'b0, 1'b0, 2'b01, 8'b10010010, 10'b0100111101, 2'b01}, // D18.4 (RD = -1) WRONG RDF
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0100111110, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0100111111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0101000000, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0101000001, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0101000010, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0101000011, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0101000100, 2'bxx}, // ?
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b01011111, 10'b0101000101, 2'b11}, // D31.2 (RD = +1)
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b11011111, 10'b0101000110, 2'b11}, // D31.6 (RD = +1)
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0101000111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0101001000, 2'bxx}, // ?
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b00111111, 10'b0101001001, 2'b11}, // D31.1 (RD = +1)
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b10111111, 10'b0101001010, 2'b11}, // D31.5 (RD = +1)
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b00011111, 10'b0101001011, 2'b01}, // D31.0 (RD = +1)
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b01111111, 10'b0101001100, 2'b11}, // D31.3 (RD = +1)
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b10011111, 10'b0101001101, 2'b01}, // D31.4 (RD = +1)
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b11111111, 10'b0101001110, 2'b01}, // D31.7 (RD = +1)
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0101001111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0101010000, 2'bxx}, // ?
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b11101010, 10'b0101010001, 2'b11}, // D10.7 (RD = +1)
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b10001010, 10'b0101010010, 2'b11}, // D10.4 (RD = +1)
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b01101010, 10'b0101010011, 2'b01}, // D10.3 (RD = +1)
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b00001010, 10'b0101010100, 2'b11}, // D10.0 (RD = +1)
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b01001010, 10'b0101010101, 2'b01}, // D10.2 (RD = +1)
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b11001010, 10'b0101010110, 2'b01}, // D10.6 (RD = +1)
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0101010111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0101011000, 2'bxx}, // ?
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b00101010, 10'b0101011001, 2'b01}, // D10.1 (RD = +1)
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b10101010, 10'b0101011010, 2'b01}, // D10.5 (RD = +1)
    {1'b1, 1'b0, 1'b0, 2'b01, 8'b00001010, 10'b0101011011, 2'b01}, // D10.0 (RD = -1) WRONG RDF
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0101011100, 2'bxx}, // ?
    {1'b1, 1'b0, 1'b0, 2'b01, 8'b10001010, 10'b0101011101, 2'b01}, // D10.4 (RD = -1) WRONG RDF
    {1'b1, 1'b0, 1'b0, 2'b01, 8'b11101010, 10'b0101011110, 2'b01}, // D10.7 (RD = -1) WRONG RDF
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0101011111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0101100000, 2'bxx}, // ?
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b11111010, 10'b0101100001, 2'b11}, // D26.7 (RD = +1)
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b10011010, 10'b0101100010, 2'b11}, // D26.4 (RD = +1)
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b01111010, 10'b0101100011, 2'b01}, // D26.3 (RD = +1)
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b00011010, 10'b0101100100, 2'b11}, // D26.0 (RD = +1)
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b01011010, 10'b0101100101, 2'b01}, // D26.2 (RD = +1)
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b11011010, 10'b0101100110, 2'b01}, // D26.6 (RD = +1)
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0101100111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0101101000, 2'bxx}, // ?
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b00111010, 10'b0101101001, 2'b01}, // D26.1 (RD = +1)
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b10111010, 10'b0101101010, 2'b01}, // D26.5 (RD = +1)
    {1'b1, 1'b0, 1'b0, 2'b01, 8'b00011010, 10'b0101101011, 2'b01}, // D26.0 (RD = -1) WRONG RDF
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0101101100, 2'bxx}, // ?
    {1'b1, 1'b0, 1'b0, 2'b01, 8'b10011010, 10'b0101101101, 2'b01}, // D26.4 (RD = -1) WRONG RDF
    {1'b1, 1'b0, 1'b0, 2'b01, 8'b11111010, 10'b0101101110, 2'b01}, // D26.7 (RD = -1) WRONG RDF
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0101101111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0101110000, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0101110001, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0101110010, 2'bxx}, // ?
    {1'b1, 1'b0, 1'b0, 2'b01, 8'b01101111, 10'b0101110011, 2'b01}, // D15.3 (RD = -1) WRONG RDF
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0101110100, 2'bxx}, // ?
    {1'b1, 1'b0, 1'b0, 2'b01, 8'b01001111, 10'b0101110101, 2'b01}, // D15.2 (RD = -1) WRONG RDF
    {1'b1, 1'b0, 1'b0, 2'b01, 8'b11001111, 10'b0101110110, 2'b01}, // D15.6 (RD = -1) WRONG RDF
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0101110111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0101111000, 2'bxx}, // ?
    {1'b1, 1'b0, 1'b0, 2'b01, 8'b00101111, 10'b0101111001, 2'b01}, // D15.1 (RD = -1) WRONG RDF
    {1'b1, 1'b0, 1'b0, 2'b01, 8'b10101111, 10'b0101111010, 2'b01}, // D15.5 (RD = -1) WRONG RDF
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0101111011, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0101111100, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0101111101, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0101111110, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0101111111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0110000000, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0110000001, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0110000010, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0110000011, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0110000100, 2'bxx}, // ?
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b01000000, 10'b0110000101, 2'b11}, // D00.2 (RD = +1)
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b11000000, 10'b0110000110, 2'b11}, // D00.6 (RD = +1)
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0110000111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0110001000, 2'bxx}, // ?
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b00100000, 10'b0110001001, 2'b11}, // D00.1 (RD = +1)
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b10100000, 10'b0110001010, 2'b11}, // D00.5 (RD = +1)
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b00000000, 10'b0110001011, 2'b01}, // D00.0 (RD = +1)
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b01100000, 10'b0110001100, 2'b11}, // D00.3 (RD = +1)
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b10000000, 10'b0110001101, 2'b01}, // D00.4 (RD = +1)
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b11100000, 10'b0110001110, 2'b01}, // D00.7 (RD = +1)
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0110001111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0110010000, 2'bxx}, // ?
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b11100110, 10'b0110010001, 2'b11}, // D06.7 (RD = +1)
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b10000110, 10'b0110010010, 2'b11}, // D06.4 (RD = +1)
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b01100110, 10'b0110010011, 2'b01}, // D06.3 (RD = +1)
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b00000110, 10'b0110010100, 2'b11}, // D06.0 (RD = +1)
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b01000110, 10'b0110010101, 2'b01}, // D06.2 (RD = +1)
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b11000110, 10'b0110010110, 2'b01}, // D06.6 (RD = +1)
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0110010111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0110011000, 2'bxx}, // ?
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b00100110, 10'b0110011001, 2'b01}, // D06.1 (RD = +1)
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b10100110, 10'b0110011010, 2'b01}, // D06.5 (RD = +1)
    {1'b1, 1'b0, 1'b0, 2'b01, 8'b00000110, 10'b0110011011, 2'b01}, // D06.0 (RD = -1) WRONG RDF
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0110011100, 2'bxx}, // ?
    {1'b1, 1'b0, 1'b0, 2'b01, 8'b10000110, 10'b0110011101, 2'b01}, // D06.4 (RD = -1) WRONG RDF
    {1'b1, 1'b0, 1'b0, 2'b01, 8'b11100110, 10'b0110011110, 2'b01}, // D06.7 (RD = -1) WRONG RDF
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0110011111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0110100000, 2'bxx}, // ?
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b11110110, 10'b0110100001, 2'b11}, // D22.7 (RD = +1)
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b10010110, 10'b0110100010, 2'b11}, // D22.4 (RD = +1)
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b01110110, 10'b0110100011, 2'b01}, // D22.3 (RD = +1)
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b00010110, 10'b0110100100, 2'b11}, // D22.0 (RD = +1)
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b01010110, 10'b0110100101, 2'b01}, // D22.2 (RD = +1)
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b11010110, 10'b0110100110, 2'b01}, // D22.6 (RD = +1)
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0110100111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0110101000, 2'bxx}, // ?
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b00110110, 10'b0110101001, 2'b01}, // D22.1 (RD = +1)
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b10110110, 10'b0110101010, 2'b01}, // D22.5 (RD = +1)
    {1'b1, 1'b0, 1'b0, 2'b01, 8'b00010110, 10'b0110101011, 2'b01}, // D22.0 (RD = -1) WRONG RDF
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0110101100, 2'bxx}, // ?
    {1'b1, 1'b0, 1'b0, 2'b01, 8'b10010110, 10'b0110101101, 2'b01}, // D22.4 (RD = -1) WRONG RDF
    {1'b1, 1'b0, 1'b0, 2'b01, 8'b11110110, 10'b0110101110, 2'b01}, // D22.7 (RD = -1) WRONG RDF
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0110101111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0110110000, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0110110001, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0110110010, 2'bxx}, // ?
    {1'b1, 1'b0, 1'b0, 2'b01, 8'b01110000, 10'b0110110011, 2'b01}, // D16.3 (RD = -1) WRONG RDF
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0110110100, 2'bxx}, // ?
    {1'b1, 1'b0, 1'b0, 2'b01, 8'b01010000, 10'b0110110101, 2'b01}, // D16.2 (RD = -1) WRONG RDF
    {1'b1, 1'b0, 1'b0, 2'b01, 8'b11010000, 10'b0110110110, 2'b01}, // D16.6 (RD = -1) WRONG RDF
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0110110111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0110111000, 2'bxx}, // ?
    {1'b1, 1'b0, 1'b0, 2'b01, 8'b00110000, 10'b0110111001, 2'b01}, // D16.1 (RD = -1) WRONG RDF
    {1'b1, 1'b0, 1'b0, 2'b01, 8'b10110000, 10'b0110111010, 2'b01}, // D16.5 (RD = -1) WRONG RDF
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0110111011, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0110111100, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0110111101, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0110111110, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0110111111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0111000000, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0111000001, 2'bxx}, // ?
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b10001110, 10'b0111000010, 2'b11}, // D14.4 (RD = +1)
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b01101110, 10'b0111000011, 2'b01}, // D14.3 (RD = +1)
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b00001110, 10'b0111000100, 2'b11}, // D14.0 (RD = +1)
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b01001110, 10'b0111000101, 2'b01}, // D14.2 (RD = +1)
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b11001110, 10'b0111000110, 2'b01}, // D14.6 (RD = +1)
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0111000111, 2'bxx}, // ?
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b11101110, 10'b0111001000, 2'b11}, // D14.7 (RD = +1)
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b00101110, 10'b0111001001, 2'b01}, // D14.1 (RD = +1)
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b10101110, 10'b0111001010, 2'b01}, // D14.5 (RD = +1)
    {1'b1, 1'b0, 1'b0, 2'b01, 8'b00001110, 10'b0111001011, 2'b01}, // D14.0 (RD = -1) WRONG RDF
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0111001100, 2'bxx}, // ?
    {1'b1, 1'b0, 1'b0, 2'b01, 8'b10001110, 10'b0111001101, 2'b01}, // D14.4 (RD = -1) WRONG RDF
    {1'b1, 1'b0, 1'b0, 2'b01, 8'b11101110, 10'b0111001110, 2'b01}, // D14.7 (RD = -1) WRONG RDF
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0111001111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0111010000, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0111010001, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0111010010, 2'bxx}, // ?
    {1'b1, 1'b0, 1'b0, 2'b01, 8'b01100001, 10'b0111010011, 2'b01}, // D01.3 (RD = -1) WRONG RDF
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0111010100, 2'bxx}, // ?
    {1'b1, 1'b0, 1'b0, 2'b01, 8'b01000001, 10'b0111010101, 2'b01}, // D01.2 (RD = -1) WRONG RDF
    {1'b1, 1'b0, 1'b0, 2'b01, 8'b11000001, 10'b0111010110, 2'b01}, // D01.6 (RD = -1) WRONG RDF
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0111010111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0111011000, 2'bxx}, // ?
    {1'b1, 1'b0, 1'b0, 2'b01, 8'b00100001, 10'b0111011001, 2'b01}, // D01.1 (RD = -1) WRONG RDF
    {1'b1, 1'b0, 1'b0, 2'b01, 8'b10100001, 10'b0111011010, 2'b01}, // D01.5 (RD = -1) WRONG RDF
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0111011011, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0111011100, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0111011101, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0111011110, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0111011111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0111100000, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0111100001, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0111100010, 2'bxx}, // ?
    {1'b1, 1'b0, 1'b0, 2'b01, 8'b01111110, 10'b0111100011, 2'b01}, // D30.3 (RD = -1) WRONG RDF
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0111100100, 2'bxx}, // ?
    {1'b1, 1'b0, 1'b0, 2'b01, 8'b01011110, 10'b0111100101, 2'b01}, // D30.2 (RD = -1) WRONG RDF
    {1'b1, 1'b0, 1'b0, 2'b01, 8'b11011110, 10'b0111100110, 2'b01}, // D30.6 (RD = -1) WRONG RDF
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0111100111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0111101000, 2'bxx}, // ?
    {1'b1, 1'b0, 1'b0, 2'b01, 8'b00111110, 10'b0111101001, 2'b01}, // D30.1 (RD = -1) WRONG RDF
    {1'b1, 1'b0, 1'b0, 2'b01, 8'b10111110, 10'b0111101010, 2'b01}, // D30.5 (RD = -1) WRONG RDF
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0111101011, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0111101100, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0111101101, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0111101110, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0111101111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0111110000, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0111110001, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0111110010, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0111110011, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0111110100, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0111110101, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0111110110, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0111110111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0111111000, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0111111001, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0111111010, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0111111011, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0111111100, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0111111101, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0111111110, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b0111111111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1000000000, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1000000001, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1000000010, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1000000011, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1000000100, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1000000101, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1000000110, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1000000111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1000001000, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1000001001, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1000001010, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1000001011, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1000001100, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1000001101, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1000001110, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1000001111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1000010000, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1000010001, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1000010010, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1000010011, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1000010100, 2'bxx}, // ?
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b01011110, 10'b1000010101, 2'b11}, // D30.2 (RD = +1)
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b11011110, 10'b1000010110, 2'b11}, // D30.6 (RD = +1)
    {1'b0, 1'b0, 1'b1, 2'b01, 8'b11111110, 10'b1000010111, 2'b01}, // K30.7 (RD = +1)
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1000011000, 2'bxx}, // ?
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b00111110, 10'b1000011001, 2'b11}, // D30.1 (RD = +1)
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b10111110, 10'b1000011010, 2'b11}, // D30.5 (RD = +1)
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b00011110, 10'b1000011011, 2'b01}, // D30.0 (RD = +1)
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b01111110, 10'b1000011100, 2'b11}, // D30.3 (RD = +1)
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b10011110, 10'b1000011101, 2'b01}, // D30.4 (RD = +1)
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b11111110, 10'b1000011110, 2'b01}, // D30.7 (RD = +1)
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1000011111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1000100000, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1000100001, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1000100010, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1000100011, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1000100100, 2'bxx}, // ?
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b01000001, 10'b1000100101, 2'b11}, // D01.2 (RD = +1)
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b11000001, 10'b1000100110, 2'b11}, // D01.6 (RD = +1)
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1000100111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1000101000, 2'bxx}, // ?
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b00100001, 10'b1000101001, 2'b11}, // D01.1 (RD = +1)
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b10100001, 10'b1000101010, 2'b11}, // D01.5 (RD = +1)
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b00000001, 10'b1000101011, 2'b01}, // D01.0 (RD = +1)
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b01100001, 10'b1000101100, 2'b11}, // D01.3 (RD = +1)
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b10000001, 10'b1000101101, 2'b01}, // D01.4 (RD = +1)
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b11100001, 10'b1000101110, 2'b01}, // D01.7 (RD = +1)
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1000101111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1000110000, 2'bxx}, // ?
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b11110001, 10'b1000110001, 2'b11}, // D17.7 (RD = +1)
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b10010001, 10'b1000110010, 2'b11}, // D17.4 (RD = +1)
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b01110001, 10'b1000110011, 2'b01}, // D17.3 (RD = +1)
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b00010001, 10'b1000110100, 2'b11}, // D17.0 (RD = +1)
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b01010001, 10'b1000110101, 2'b01}, // D17.2 (RD = +1)
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b11010001, 10'b1000110110, 2'b01}, // D17.6 (RD = +1)
    {1'b1, 1'b0, 1'b0, 2'b01, 8'b11110001, 10'b1000110111, 2'b01}, // D17.7 (RD = -1) WRONG RDF
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1000111000, 2'bxx}, // ?
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b00110001, 10'b1000111001, 2'b01}, // D17.1 (RD = +1)
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b10110001, 10'b1000111010, 2'b01}, // D17.5 (RD = +1)
    {1'b1, 1'b0, 1'b0, 2'b01, 8'b00010001, 10'b1000111011, 2'b01}, // D17.0 (RD = -1) WRONG RDF
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1000111100, 2'bxx}, // ?
    {1'b1, 1'b0, 1'b0, 2'b01, 8'b10010001, 10'b1000111101, 2'b01}, // D17.4 (RD = -1) WRONG RDF
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1000111110, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1000111111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1001000000, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1001000001, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1001000010, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1001000011, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1001000100, 2'bxx}, // ?
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b01010000, 10'b1001000101, 2'b11}, // D16.2 (RD = +1)
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b11010000, 10'b1001000110, 2'b11}, // D16.6 (RD = +1)
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1001000111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1001001000, 2'bxx}, // ?
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b00110000, 10'b1001001001, 2'b11}, // D16.1 (RD = +1)
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b10110000, 10'b1001001010, 2'b11}, // D16.5 (RD = +1)
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b00010000, 10'b1001001011, 2'b01}, // D16.0 (RD = +1)
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b01110000, 10'b1001001100, 2'b11}, // D16.3 (RD = +1)
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b10010000, 10'b1001001101, 2'b01}, // D16.4 (RD = +1)
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b11110000, 10'b1001001110, 2'b01}, // D16.7 (RD = +1)
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1001001111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1001010000, 2'bxx}, // ?
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b11101001, 10'b1001010001, 2'b11}, // D09.7 (RD = +1)
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b10001001, 10'b1001010010, 2'b11}, // D09.4 (RD = +1)
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b01101001, 10'b1001010011, 2'b01}, // D09.3 (RD = +1)
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b00001001, 10'b1001010100, 2'b11}, // D09.0 (RD = +1)
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b01001001, 10'b1001010101, 2'b01}, // D09.2 (RD = +1)
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b11001001, 10'b1001010110, 2'b01}, // D09.6 (RD = +1)
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1001010111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1001011000, 2'bxx}, // ?
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b00101001, 10'b1001011001, 2'b01}, // D09.1 (RD = +1)
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b10101001, 10'b1001011010, 2'b01}, // D09.5 (RD = +1)
    {1'b1, 1'b0, 1'b0, 2'b01, 8'b00001001, 10'b1001011011, 2'b01}, // D09.0 (RD = -1) WRONG RDF
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1001011100, 2'bxx}, // ?
    {1'b1, 1'b0, 1'b0, 2'b01, 8'b10001001, 10'b1001011101, 2'b01}, // D09.4 (RD = -1) WRONG RDF
    {1'b1, 1'b0, 1'b0, 2'b01, 8'b11101001, 10'b1001011110, 2'b01}, // D09.7 (RD = -1) WRONG RDF
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1001011111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1001100000, 2'bxx}, // ?
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b11111001, 10'b1001100001, 2'b11}, // D25.7 (RD = +1)
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b10011001, 10'b1001100010, 2'b11}, // D25.4 (RD = +1)
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b01111001, 10'b1001100011, 2'b01}, // D25.3 (RD = +1)
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b00011001, 10'b1001100100, 2'b11}, // D25.0 (RD = +1)
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b01011001, 10'b1001100101, 2'b01}, // D25.2 (RD = +1)
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b11011001, 10'b1001100110, 2'b01}, // D25.6 (RD = +1)
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1001100111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1001101000, 2'bxx}, // ?
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b00111001, 10'b1001101001, 2'b01}, // D25.1 (RD = +1)
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b10111001, 10'b1001101010, 2'b01}, // D25.5 (RD = +1)
    {1'b1, 1'b0, 1'b0, 2'b01, 8'b00011001, 10'b1001101011, 2'b01}, // D25.0 (RD = -1) WRONG RDF
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1001101100, 2'bxx}, // ?
    {1'b1, 1'b0, 1'b0, 2'b01, 8'b10011001, 10'b1001101101, 2'b01}, // D25.4 (RD = -1) WRONG RDF
    {1'b1, 1'b0, 1'b0, 2'b01, 8'b11111001, 10'b1001101110, 2'b01}, // D25.7 (RD = -1) WRONG RDF
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1001101111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1001110000, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1001110001, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1001110010, 2'bxx}, // ?
    {1'b1, 1'b0, 1'b0, 2'b01, 8'b01100000, 10'b1001110011, 2'b01}, // D00.3 (RD = -1) WRONG RDF
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1001110100, 2'bxx}, // ?
    {1'b1, 1'b0, 1'b0, 2'b01, 8'b01000000, 10'b1001110101, 2'b01}, // D00.2 (RD = -1) WRONG RDF
    {1'b1, 1'b0, 1'b0, 2'b01, 8'b11000000, 10'b1001110110, 2'b01}, // D00.6 (RD = -1) WRONG RDF
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1001110111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1001111000, 2'bxx}, // ?
    {1'b1, 1'b0, 1'b0, 2'b01, 8'b00100000, 10'b1001111001, 2'b01}, // D00.1 (RD = -1) WRONG RDF
    {1'b1, 1'b0, 1'b0, 2'b01, 8'b10100000, 10'b1001111010, 2'b01}, // D00.5 (RD = -1) WRONG RDF
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1001111011, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1001111100, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1001111101, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1001111110, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1001111111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1010000000, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1010000001, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1010000010, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1010000011, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1010000100, 2'bxx}, // ?
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b01001111, 10'b1010000101, 2'b11}, // D15.2 (RD = +1)
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b11001111, 10'b1010000110, 2'b11}, // D15.6 (RD = +1)
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1010000111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1010001000, 2'bxx}, // ?
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b00101111, 10'b1010001001, 2'b11}, // D15.1 (RD = +1)
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b10101111, 10'b1010001010, 2'b11}, // D15.5 (RD = +1)
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b00001111, 10'b1010001011, 2'b01}, // D15.0 (RD = +1)
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b01101111, 10'b1010001100, 2'b11}, // D15.3 (RD = +1)
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b10001111, 10'b1010001101, 2'b01}, // D15.4 (RD = +1)
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b11101111, 10'b1010001110, 2'b01}, // D15.7 (RD = +1)
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1010001111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1010010000, 2'bxx}, // ?
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b11100101, 10'b1010010001, 2'b11}, // D05.7 (RD = +1)
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b10000101, 10'b1010010010, 2'b11}, // D05.4 (RD = +1)
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b01100101, 10'b1010010011, 2'b01}, // D05.3 (RD = +1)
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b00000101, 10'b1010010100, 2'b11}, // D05.0 (RD = +1)
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b01000101, 10'b1010010101, 2'b01}, // D05.2 (RD = +1)
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b11000101, 10'b1010010110, 2'b01}, // D05.6 (RD = +1)
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1010010111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1010011000, 2'bxx}, // ?
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b00100101, 10'b1010011001, 2'b01}, // D05.1 (RD = +1)
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b10100101, 10'b1010011010, 2'b01}, // D05.5 (RD = +1)
    {1'b1, 1'b0, 1'b0, 2'b01, 8'b00000101, 10'b1010011011, 2'b01}, // D05.0 (RD = -1) WRONG RDF
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1010011100, 2'bxx}, // ?
    {1'b1, 1'b0, 1'b0, 2'b01, 8'b10000101, 10'b1010011101, 2'b01}, // D05.4 (RD = -1) WRONG RDF
    {1'b1, 1'b0, 1'b0, 2'b01, 8'b11100101, 10'b1010011110, 2'b01}, // D05.7 (RD = -1) WRONG RDF
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1010011111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1010100000, 2'bxx}, // ?
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b11110101, 10'b1010100001, 2'b11}, // D21.7 (RD = +1)
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b10010101, 10'b1010100010, 2'b11}, // D21.4 (RD = +1)
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b01110101, 10'b1010100011, 2'b01}, // D21.3 (RD = +1)
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b00010101, 10'b1010100100, 2'b11}, // D21.0 (RD = +1)
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b01010101, 10'b1010100101, 2'b01}, // D21.2 (RD = +1)
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b11010101, 10'b1010100110, 2'b01}, // D21.6 (RD = +1)
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1010100111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1010101000, 2'bxx}, // ?
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b00110101, 10'b1010101001, 2'b01}, // D21.1 (RD = +1)
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b10110101, 10'b1010101010, 2'b01}, // D21.5 (RD = +1)
    {1'b1, 1'b0, 1'b0, 2'b01, 8'b00010101, 10'b1010101011, 2'b01}, // D21.0 (RD = -1) WRONG RDF
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1010101100, 2'bxx}, // ?
    {1'b1, 1'b0, 1'b0, 2'b01, 8'b10010101, 10'b1010101101, 2'b01}, // D21.4 (RD = -1) WRONG RDF
    {1'b1, 1'b0, 1'b0, 2'b01, 8'b11110101, 10'b1010101110, 2'b01}, // D21.7 (RD = -1) WRONG RDF
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1010101111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1010110000, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1010110001, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1010110010, 2'bxx}, // ?
    {1'b1, 1'b0, 1'b0, 2'b01, 8'b01111111, 10'b1010110011, 2'b01}, // D31.3 (RD = -1) WRONG RDF
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1010110100, 2'bxx}, // ?
    {1'b1, 1'b0, 1'b0, 2'b01, 8'b01011111, 10'b1010110101, 2'b01}, // D31.2 (RD = -1) WRONG RDF
    {1'b1, 1'b0, 1'b0, 2'b01, 8'b11011111, 10'b1010110110, 2'b01}, // D31.6 (RD = -1) WRONG RDF
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1010110111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1010111000, 2'bxx}, // ?
    {1'b1, 1'b0, 1'b0, 2'b01, 8'b00111111, 10'b1010111001, 2'b01}, // D31.1 (RD = -1) WRONG RDF
    {1'b1, 1'b0, 1'b0, 2'b01, 8'b10111111, 10'b1010111010, 2'b01}, // D31.5 (RD = -1) WRONG RDF
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1010111011, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1010111100, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1010111101, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1010111110, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1010111111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1011000000, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1011000001, 2'bxx}, // ?
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b10001101, 10'b1011000010, 2'b11}, // D13.4 (RD = +1)
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b01101101, 10'b1011000011, 2'b01}, // D13.3 (RD = +1)
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b00001101, 10'b1011000100, 2'b11}, // D13.0 (RD = +1)
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b01001101, 10'b1011000101, 2'b01}, // D13.2 (RD = +1)
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b11001101, 10'b1011000110, 2'b01}, // D13.6 (RD = +1)
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1011000111, 2'bxx}, // ?
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b11101101, 10'b1011001000, 2'b11}, // D13.7 (RD = +1)
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b00101101, 10'b1011001001, 2'b01}, // D13.1 (RD = +1)
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b10101101, 10'b1011001010, 2'b01}, // D13.5 (RD = +1)
    {1'b1, 1'b0, 1'b0, 2'b01, 8'b00001101, 10'b1011001011, 2'b01}, // D13.0 (RD = -1) WRONG RDF
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1011001100, 2'bxx}, // ?
    {1'b1, 1'b0, 1'b0, 2'b01, 8'b10001101, 10'b1011001101, 2'b01}, // D13.4 (RD = -1) WRONG RDF
    {1'b1, 1'b0, 1'b0, 2'b01, 8'b11101101, 10'b1011001110, 2'b01}, // D13.7 (RD = -1) WRONG RDF
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1011001111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1011010000, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1011010001, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1011010010, 2'bxx}, // ?
    {1'b1, 1'b0, 1'b0, 2'b01, 8'b01100010, 10'b1011010011, 2'b01}, // D02.3 (RD = -1) WRONG RDF
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1011010100, 2'bxx}, // ?
    {1'b1, 1'b0, 1'b0, 2'b01, 8'b01000010, 10'b1011010101, 2'b01}, // D02.2 (RD = -1) WRONG RDF
    {1'b1, 1'b0, 1'b0, 2'b01, 8'b11000010, 10'b1011010110, 2'b01}, // D02.6 (RD = -1) WRONG RDF
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1011010111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1011011000, 2'bxx}, // ?
    {1'b1, 1'b0, 1'b0, 2'b01, 8'b00100010, 10'b1011011001, 2'b01}, // D02.1 (RD = -1) WRONG RDF
    {1'b1, 1'b0, 1'b0, 2'b01, 8'b10100010, 10'b1011011010, 2'b01}, // D02.5 (RD = -1) WRONG RDF
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1011011011, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1011011100, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1011011101, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1011011110, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1011011111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1011100000, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1011100001, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1011100010, 2'bxx}, // ?
    {1'b1, 1'b0, 1'b0, 2'b01, 8'b01111101, 10'b1011100011, 2'b01}, // D29.3 (RD = -1) WRONG RDF
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1011100100, 2'bxx}, // ?
    {1'b1, 1'b0, 1'b0, 2'b01, 8'b01011101, 10'b1011100101, 2'b01}, // D29.2 (RD = -1) WRONG RDF
    {1'b1, 1'b0, 1'b0, 2'b01, 8'b11011101, 10'b1011100110, 2'b01}, // D29.6 (RD = -1) WRONG RDF
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1011100111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1011101000, 2'bxx}, // ?
    {1'b1, 1'b0, 1'b0, 2'b01, 8'b00111101, 10'b1011101001, 2'b01}, // D29.1 (RD = -1) WRONG RDF
    {1'b1, 1'b0, 1'b0, 2'b01, 8'b10111101, 10'b1011101010, 2'b01}, // D29.5 (RD = -1) WRONG RDF
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1011101011, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1011101100, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1011101101, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1011101110, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1011101111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1011110000, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1011110001, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1011110010, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1011110011, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1011110100, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1011110101, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1011110110, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1011110111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1011111000, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1011111001, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1011111010, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1011111011, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1011111100, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1011111101, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1011111110, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1011111111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1100000000, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1100000001, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1100000010, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1100000011, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1100000100, 2'bxx}, // ?
    {1'b0, 1'b0, 1'b1, 2'b01, 8'b10111100, 10'b1100000101, 2'b11}, // K28.5 (RD = +1)
    {1'b0, 1'b0, 1'b1, 2'b01, 8'b00111100, 10'b1100000110, 2'b11}, // K28.1 (RD = +1)
    {1'b0, 1'b0, 1'b1, 2'b01, 8'b11111100, 10'b1100000111, 2'b01}, // K28.7 (RD = +1)
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1100001000, 2'bxx}, // ?
    {1'b0, 1'b0, 1'b1, 2'b01, 8'b11011100, 10'b1100001001, 2'b11}, // K28.6 (RD = +1)
    {1'b0, 1'b0, 1'b1, 2'b01, 8'b01011100, 10'b1100001010, 2'b11}, // K28.2 (RD = +1)
    {1'b0, 1'b0, 1'b1, 2'b01, 8'b00011100, 10'b1100001011, 2'b01}, // K28.0 (RD = +1)
    {1'b0, 1'b0, 1'b1, 2'b01, 8'b01111100, 10'b1100001100, 2'b11}, // K28.3 (RD = +1)
    {1'b0, 1'b0, 1'b1, 2'b01, 8'b10011100, 10'b1100001101, 2'b01}, // K28.4 (RD = +1)
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1100001110, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1100001111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1100010000, 2'bxx}, // ?
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b11100011, 10'b1100010001, 2'b11}, // D03.7 (RD = +1)
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b10000011, 10'b1100010010, 2'b11}, // D03.4 (RD = +1)
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b01100011, 10'b1100010011, 2'b01}, // D03.3 (RD = +1)
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b00000011, 10'b1100010100, 2'b11}, // D03.0 (RD = +1)
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b01000011, 10'b1100010101, 2'b01}, // D03.2 (RD = +1)
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b11000011, 10'b1100010110, 2'b01}, // D03.6 (RD = +1)
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1100010111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1100011000, 2'bxx}, // ?
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b00100011, 10'b1100011001, 2'b01}, // D03.1 (RD = +1)
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b10100011, 10'b1100011010, 2'b01}, // D03.5 (RD = +1)
    {1'b1, 1'b0, 1'b0, 2'b01, 8'b00000011, 10'b1100011011, 2'b01}, // D03.0 (RD = -1) WRONG RDF
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1100011100, 2'bxx}, // ?
    {1'b1, 1'b0, 1'b0, 2'b01, 8'b10000011, 10'b1100011101, 2'b01}, // D03.4 (RD = -1) WRONG RDF
    {1'b1, 1'b0, 1'b0, 2'b01, 8'b11100011, 10'b1100011110, 2'b01}, // D03.7 (RD = -1) WRONG RDF
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1100011111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1100100000, 2'bxx}, // ?
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b11110011, 10'b1100100001, 2'b11}, // D19.7 (RD = +1)
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b10010011, 10'b1100100010, 2'b11}, // D19.4 (RD = +1)
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b01110011, 10'b1100100011, 2'b01}, // D19.3 (RD = +1)
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b00010011, 10'b1100100100, 2'b11}, // D19.0 (RD = +1)
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b01010011, 10'b1100100101, 2'b01}, // D19.2 (RD = +1)
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b11010011, 10'b1100100110, 2'b01}, // D19.6 (RD = +1)
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1100100111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1100101000, 2'bxx}, // ?
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b00110011, 10'b1100101001, 2'b01}, // D19.1 (RD = +1)
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b10110011, 10'b1100101010, 2'b01}, // D19.5 (RD = +1)
    {1'b1, 1'b0, 1'b0, 2'b01, 8'b00010011, 10'b1100101011, 2'b01}, // D19.0 (RD = -1) WRONG RDF
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1100101100, 2'bxx}, // ?
    {1'b1, 1'b0, 1'b0, 2'b01, 8'b10010011, 10'b1100101101, 2'b01}, // D19.4 (RD = -1) WRONG RDF
    {1'b1, 1'b0, 1'b0, 2'b01, 8'b11110011, 10'b1100101110, 2'b01}, // D19.7 (RD = -1) WRONG RDF
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1100101111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1100110000, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1100110001, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1100110010, 2'bxx}, // ?
    {1'b1, 1'b0, 1'b0, 2'b01, 8'b01111000, 10'b1100110011, 2'b01}, // D24.3 (RD = -1) WRONG RDF
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1100110100, 2'bxx}, // ?
    {1'b1, 1'b0, 1'b0, 2'b01, 8'b01011000, 10'b1100110101, 2'b01}, // D24.2 (RD = -1) WRONG RDF
    {1'b1, 1'b0, 1'b0, 2'b01, 8'b11011000, 10'b1100110110, 2'b01}, // D24.6 (RD = -1) WRONG RDF
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1100110111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1100111000, 2'bxx}, // ?
    {1'b1, 1'b0, 1'b0, 2'b01, 8'b00111000, 10'b1100111001, 2'b01}, // D24.1 (RD = -1) WRONG RDF
    {1'b1, 1'b0, 1'b0, 2'b01, 8'b10111000, 10'b1100111010, 2'b01}, // D24.5 (RD = -1) WRONG RDF
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1100111011, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1100111100, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1100111101, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1100111110, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1100111111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1101000000, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1101000001, 2'bxx}, // ?
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b10001011, 10'b1101000010, 2'b11}, // D11.4 (RD = +1)
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b01101011, 10'b1101000011, 2'b01}, // D11.3 (RD = +1)
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b00001011, 10'b1101000100, 2'b11}, // D11.0 (RD = +1)
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b01001011, 10'b1101000101, 2'b01}, // D11.2 (RD = +1)
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b11001011, 10'b1101000110, 2'b01}, // D11.6 (RD = +1)
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1101000111, 2'bxx}, // ?
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b11101011, 10'b1101001000, 2'b11}, // D11.7 (RD = +1)
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b00101011, 10'b1101001001, 2'b01}, // D11.1 (RD = +1)
    {1'b0, 1'b0, 1'b0, 2'b01, 8'b10101011, 10'b1101001010, 2'b01}, // D11.5 (RD = +1)
    {1'b1, 1'b0, 1'b0, 2'b01, 8'b00001011, 10'b1101001011, 2'b01}, // D11.0 (RD = -1) WRONG RDF
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1101001100, 2'bxx}, // ?
    {1'b1, 1'b0, 1'b0, 2'b01, 8'b10001011, 10'b1101001101, 2'b01}, // D11.4 (RD = -1) WRONG RDF
    {1'b1, 1'b0, 1'b0, 2'b01, 8'b11101011, 10'b1101001110, 2'b01}, // D11.7 (RD = -1) WRONG RDF
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1101001111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1101010000, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1101010001, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1101010010, 2'bxx}, // ?
    {1'b1, 1'b0, 1'b0, 2'b01, 8'b01100100, 10'b1101010011, 2'b01}, // D04.3 (RD = -1) WRONG RDF
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1101010100, 2'bxx}, // ?
    {1'b1, 1'b0, 1'b0, 2'b01, 8'b01000100, 10'b1101010101, 2'b01}, // D04.2 (RD = -1) WRONG RDF
    {1'b1, 1'b0, 1'b0, 2'b01, 8'b11000100, 10'b1101010110, 2'b01}, // D04.6 (RD = -1) WRONG RDF
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1101010111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1101011000, 2'bxx}, // ?
    {1'b1, 1'b0, 1'b0, 2'b01, 8'b00100100, 10'b1101011001, 2'b01}, // D04.1 (RD = -1) WRONG RDF
    {1'b1, 1'b0, 1'b0, 2'b01, 8'b10100100, 10'b1101011010, 2'b01}, // D04.5 (RD = -1) WRONG RDF
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1101011011, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1101011100, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1101011101, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1101011110, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1101011111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1101100000, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1101100001, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1101100010, 2'bxx}, // ?
    {1'b1, 1'b0, 1'b0, 2'b01, 8'b01111011, 10'b1101100011, 2'b01}, // D27.3 (RD = -1) WRONG RDF
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1101100100, 2'bxx}, // ?
    {1'b1, 1'b0, 1'b0, 2'b01, 8'b01011011, 10'b1101100101, 2'b01}, // D27.2 (RD = -1) WRONG RDF
    {1'b1, 1'b0, 1'b0, 2'b01, 8'b11011011, 10'b1101100110, 2'b01}, // D27.6 (RD = -1) WRONG RDF
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1101100111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1101101000, 2'bxx}, // ?
    {1'b1, 1'b0, 1'b0, 2'b01, 8'b00111011, 10'b1101101001, 2'b01}, // D27.1 (RD = -1) WRONG RDF
    {1'b1, 1'b0, 1'b0, 2'b01, 8'b10111011, 10'b1101101010, 2'b01}, // D27.5 (RD = -1) WRONG RDF
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1101101011, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1101101100, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1101101101, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1101101110, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1101101111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1101110000, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1101110001, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1101110010, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1101110011, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1101110100, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1101110101, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1101110110, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1101110111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1101111000, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1101111001, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1101111010, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1101111011, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1101111100, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1101111101, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1101111110, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1101111111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1110000000, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1110000001, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1110000010, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1110000011, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1110000100, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1110000101, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1110000110, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1110000111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1110001000, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1110001001, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1110001010, 2'bxx}, // ?
    {1'b1, 1'b0, 1'b0, 2'b01, 8'b00000111, 10'b1110001011, 2'b01}, // D07.0 (RD = -1) WRONG RDF
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1110001100, 2'bxx}, // ?
    {1'b1, 1'b0, 1'b0, 2'b01, 8'b10000111, 10'b1110001101, 2'b01}, // D07.4 (RD = -1) WRONG RDF
    {1'b1, 1'b0, 1'b0, 2'b01, 8'b11100111, 10'b1110001110, 2'b01}, // D07.7 (RD = -1) WRONG RDF
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1110001111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1110010000, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1110010001, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1110010010, 2'bxx}, // ?
    {1'b1, 1'b0, 1'b0, 2'b01, 8'b01101000, 10'b1110010011, 2'b01}, // D08.3 (RD = -1) WRONG RDF
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1110010100, 2'bxx}, // ?
    {1'b1, 1'b0, 1'b0, 2'b01, 8'b01001000, 10'b1110010101, 2'b01}, // D08.2 (RD = -1) WRONG RDF
    {1'b1, 1'b0, 1'b0, 2'b01, 8'b11001000, 10'b1110010110, 2'b01}, // D08.6 (RD = -1) WRONG RDF
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1110010111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1110011000, 2'bxx}, // ?
    {1'b1, 1'b0, 1'b0, 2'b01, 8'b00101000, 10'b1110011001, 2'b01}, // D08.1 (RD = -1) WRONG RDF
    {1'b1, 1'b0, 1'b0, 2'b01, 8'b10101000, 10'b1110011010, 2'b01}, // D08.5 (RD = -1) WRONG RDF
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1110011011, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1110011100, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1110011101, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1110011110, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1110011111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1110100000, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1110100001, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1110100010, 2'bxx}, // ?
    {1'b1, 1'b0, 1'b0, 2'b01, 8'b01110111, 10'b1110100011, 2'b01}, // D23.3 (RD = -1) WRONG RDF
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1110100100, 2'bxx}, // ?
    {1'b1, 1'b0, 1'b0, 2'b01, 8'b01010111, 10'b1110100101, 2'b01}, // D23.2 (RD = -1) WRONG RDF
    {1'b1, 1'b0, 1'b0, 2'b01, 8'b11010111, 10'b1110100110, 2'b01}, // D23.6 (RD = -1) WRONG RDF
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1110100111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1110101000, 2'bxx}, // ?
    {1'b1, 1'b0, 1'b0, 2'b01, 8'b00110111, 10'b1110101001, 2'b01}, // D23.1 (RD = -1) WRONG RDF
    {1'b1, 1'b0, 1'b0, 2'b01, 8'b10110111, 10'b1110101010, 2'b01}, // D23.5 (RD = -1) WRONG RDF
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1110101011, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1110101100, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1110101101, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1110101110, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1110101111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1110110000, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1110110001, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1110110010, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1110110011, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1110110100, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1110110101, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1110110110, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1110110111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1110111000, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1110111001, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1110111010, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1110111011, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1110111100, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1110111101, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1110111110, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1110111111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1111000000, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1111000001, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1111000010, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1111000011, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1111000100, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1111000101, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1111000110, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1111000111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1111001000, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1111001001, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1111001010, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1111001011, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1111001100, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1111001101, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1111001110, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1111001111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1111010000, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1111010001, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1111010010, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1111010011, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1111010100, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1111010101, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1111010110, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1111010111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1111011000, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1111011001, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1111011010, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1111011011, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1111011100, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1111011101, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1111011110, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1111011111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1111100000, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1111100001, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1111100010, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1111100011, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1111100100, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1111100101, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1111100110, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1111100111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1111101000, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1111101001, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1111101010, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1111101011, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1111101100, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1111101101, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1111101110, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1111101111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1111110000, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1111110001, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1111110010, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1111110011, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1111110100, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1111110101, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1111110110, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1111110111, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1111111000, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1111111001, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1111111010, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1111111011, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1111111100, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1111111101, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1111111110, 2'bxx}, // ?
    {1'bx, 1'b1, 1'bx, 2'b01, 8'bxxxxxxxx, 10'b1111111111, 2'bxx}  // ?
  };

  string dec_byte_name [2048] = '{
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "D23.2 (RD = +1) WRONG RDF",
    "D23.6 (RD = +1) WRONG RDF",
    "?",
    "?",
    "D23.1 (RD = +1) WRONG RDF",
    "D23.5 (RD = +1) WRONG RDF",
    "?",
    "D23.3 (RD = +1) WRONG RDF",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "D08.2 (RD = +1) WRONG RDF",
    "D08.6 (RD = +1) WRONG RDF",
    "?",
    "?",
    "D08.1 (RD = +1) WRONG RDF",
    "D08.5 (RD = +1) WRONG RDF",
    "?",
    "D08.3 (RD = +1) WRONG RDF",
    "?",
    "?",
    "?",
    "?",
    "D07.7 (RD = +1) WRONG RDF",
    "D07.4 (RD = +1) WRONG RDF",
    "?",
    "D07.0 (RD = +1) WRONG RDF",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "D27.2 (RD = +1) WRONG RDF",
    "D27.6 (RD = +1) WRONG RDF",
    "?",
    "?",
    "D27.1 (RD = +1) WRONG RDF",
    "D27.5 (RD = +1) WRONG RDF",
    "?",
    "D27.3 (RD = +1) WRONG RDF",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "D04.2 (RD = +1) WRONG RDF",
    "D04.6 (RD = +1) WRONG RDF",
    "?",
    "?",
    "D04.1 (RD = +1) WRONG RDF",
    "D04.5 (RD = +1) WRONG RDF",
    "?",
    "D04.3 (RD = +1) WRONG RDF",
    "?",
    "?",
    "?",
    "?",
    "D20.7 (RD = +1) WRONG RDF",
    "D20.4 (RD = +1) WRONG RDF",
    "?",
    "D20.0 (RD = +1) WRONG RDF",
    "D20.2 (RD = -1)",
    "D20.6 (RD = -1)",
    "D20.7 (RD = -1)",
    "?",
    "D20.1 (RD = -1)",
    "D20.5 (RD = -1)",
    "D20.0 (RD = -1)",
    "D20.3 (RD = -1)",
    "D20.4 (RD = -1)",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "D24.2 (RD = +1) WRONG RDF",
    "D24.6 (RD = +1) WRONG RDF",
    "?",
    "?",
    "D24.1 (RD = +1) WRONG RDF",
    "D24.5 (RD = +1) WRONG RDF",
    "?",
    "D24.3 (RD = +1) WRONG RDF",
    "?",
    "?",
    "?",
    "?",
    "D12.7 (RD = +1) WRONG RDF",
    "D12.4 (RD = +1) WRONG RDF",
    "?",
    "D12.0 (RD = +1) WRONG RDF",
    "D12.2 (RD = -1)",
    "D12.6 (RD = -1)",
    "?",
    "?",
    "D12.1 (RD = -1)",
    "D12.5 (RD = -1)",
    "D12.0 (RD = -1)",
    "D12.3 (RD = -1)",
    "D12.4 (RD = -1)",
    "D12.7 (RD = -1)",
    "?",
    "?",
    "D28.7 (RD = +1) WRONG RDF",
    "D28.4 (RD = +1) WRONG RDF",
    "?",
    "D28.0 (RD = +1) WRONG RDF",
    "D28.2 (RD = -1)",
    "D28.6 (RD = -1)",
    "?",
    "?",
    "D28.1 (RD = -1)",
    "D28.5 (RD = -1)",
    "D28.0 (RD = -1)",
    "D28.3 (RD = -1)",
    "D28.4 (RD = -1)",
    "D28.7 (RD = -1)",
    "?",
    "?",
    "?",
    "K28.4 (RD = -1)",
    "K28.3 (RD = -1)",
    "K28.0 (RD = -1)",
    "K28.2 (RD = -1)",
    "K28.6 (RD = -1)",
    "?",
    "K28.7 (RD = -1)",
    "K28.1 (RD = -1)",
    "K28.5 (RD = -1)",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "D29.2 (RD = +1) WRONG RDF",
    "D29.6 (RD = +1) WRONG RDF",
    "?",
    "?",
    "D29.1 (RD = +1) WRONG RDF",
    "D29.5 (RD = +1) WRONG RDF",
    "?",
    "D29.3 (RD = +1) WRONG RDF",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "D02.2 (RD = +1) WRONG RDF",
    "D02.6 (RD = +1) WRONG RDF",
    "?",
    "?",
    "D02.1 (RD = +1) WRONG RDF",
    "D02.5 (RD = +1) WRONG RDF",
    "?",
    "D02.3 (RD = +1) WRONG RDF",
    "?",
    "?",
    "?",
    "?",
    "D18.7 (RD = +1) WRONG RDF",
    "D18.4 (RD = +1) WRONG RDF",
    "?",
    "D18.0 (RD = +1) WRONG RDF",
    "D18.2 (RD = -1)",
    "D18.6 (RD = -1)",
    "D18.7 (RD = -1)",
    "?",
    "D18.1 (RD = -1)",
    "D18.5 (RD = -1)",
    "D18.0 (RD = -1)",
    "D18.3 (RD = -1)",
    "D18.4 (RD = -1)",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "D31.2 (RD = +1) WRONG RDF",
    "D31.6 (RD = +1) WRONG RDF",
    "?",
    "?",
    "D31.1 (RD = +1) WRONG RDF",
    "D31.5 (RD = +1) WRONG RDF",
    "?",
    "D31.3 (RD = +1) WRONG RDF",
    "?",
    "?",
    "?",
    "?",
    "D10.7 (RD = +1) WRONG RDF",
    "D10.4 (RD = +1) WRONG RDF",
    "?",
    "D10.0 (RD = +1) WRONG RDF",
    "D10.2 (RD = -1)",
    "D10.6 (RD = -1)",
    "?",
    "?",
    "D10.1 (RD = -1)",
    "D10.5 (RD = -1)",
    "D10.0 (RD = -1)",
    "D10.3 (RD = -1)",
    "D10.4 (RD = -1)",
    "D10.7 (RD = -1)",
    "?",
    "?",
    "D26.7 (RD = +1) WRONG RDF",
    "D26.4 (RD = +1) WRONG RDF",
    "?",
    "D26.0 (RD = +1) WRONG RDF",
    "D26.2 (RD = -1)",
    "D26.6 (RD = -1)",
    "?",
    "?",
    "D26.1 (RD = -1)",
    "D26.5 (RD = -1)",
    "D26.0 (RD = -1)",
    "D26.3 (RD = -1)",
    "D26.4 (RD = -1)",
    "D26.7 (RD = -1)",
    "?",
    "?",
    "D15.7 (RD = -1)",
    "D15.4 (RD = -1)",
    "D15.3 (RD = -1)",
    "D15.0 (RD = -1)",
    "D15.2 (RD = -1)",
    "D15.6 (RD = -1)",
    "?",
    "?",
    "D15.1 (RD = -1)",
    "D15.5 (RD = -1)",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "D00.2 (RD = +1) WRONG RDF",
    "D00.6 (RD = +1) WRONG RDF",
    "?",
    "?",
    "D00.1 (RD = +1) WRONG RDF",
    "D00.5 (RD = +1) WRONG RDF",
    "?",
    "D00.3 (RD = +1) WRONG RDF",
    "?",
    "?",
    "?",
    "?",
    "D06.7 (RD = +1) WRONG RDF",
    "D06.4 (RD = +1) WRONG RDF",
    "?",
    "D06.0 (RD = +1) WRONG RDF",
    "D06.2 (RD = -1)",
    "D06.6 (RD = -1)",
    "?",
    "?",
    "D06.1 (RD = -1)",
    "D06.5 (RD = -1)",
    "D06.0 (RD = -1)",
    "D06.3 (RD = -1)",
    "D06.4 (RD = -1)",
    "D06.7 (RD = -1)",
    "?",
    "?",
    "D22.7 (RD = +1) WRONG RDF",
    "D22.4 (RD = +1) WRONG RDF",
    "?",
    "D22.0 (RD = +1) WRONG RDF",
    "D22.2 (RD = -1)",
    "D22.6 (RD = -1)",
    "?",
    "?",
    "D22.1 (RD = -1)",
    "D22.5 (RD = -1)",
    "D22.0 (RD = -1)",
    "D22.3 (RD = -1)",
    "D22.4 (RD = -1)",
    "D22.7 (RD = -1)",
    "?",
    "?",
    "D16.7 (RD = -1)",
    "D16.4 (RD = -1)",
    "D16.3 (RD = -1)",
    "D16.0 (RD = -1)",
    "D16.2 (RD = -1)",
    "D16.6 (RD = -1)",
    "?",
    "?",
    "D16.1 (RD = -1)",
    "D16.5 (RD = -1)",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "D14.4 (RD = +1) WRONG RDF",
    "?",
    "D14.0 (RD = +1) WRONG RDF",
    "D14.2 (RD = -1)",
    "D14.6 (RD = -1)",
    "?",
    "D14.7 (RD = +1) WRONG RDF",
    "D14.1 (RD = -1)",
    "D14.5 (RD = -1)",
    "D14.0 (RD = -1)",
    "D14.3 (RD = -1)",
    "D14.4 (RD = -1)",
    "D14.7 (RD = -1)",
    "?",
    "?",
    "D01.7 (RD = -1)",
    "D01.4 (RD = -1)",
    "D01.3 (RD = -1)",
    "D01.0 (RD = -1)",
    "D01.2 (RD = -1)",
    "D01.6 (RD = -1)",
    "?",
    "?",
    "D01.1 (RD = -1)",
    "D01.5 (RD = -1)",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "D30.7 (RD = -1)",
    "D30.4 (RD = -1)",
    "D30.3 (RD = -1)",
    "D30.0 (RD = -1)",
    "D30.2 (RD = -1)",
    "D30.6 (RD = -1)",
    "?",
    "K30.7 (RD = -1)",
    "D30.1 (RD = -1)",
    "D30.5 (RD = -1)",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "D30.2 (RD = +1) WRONG RDF",
    "D30.6 (RD = +1) WRONG RDF",
    "?",
    "?",
    "D30.1 (RD = +1) WRONG RDF",
    "D30.5 (RD = +1) WRONG RDF",
    "?",
    "D30.3 (RD = +1) WRONG RDF",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "D01.2 (RD = +1) WRONG RDF",
    "D01.6 (RD = +1) WRONG RDF",
    "?",
    "?",
    "D01.1 (RD = +1) WRONG RDF",
    "D01.5 (RD = +1) WRONG RDF",
    "?",
    "D01.3 (RD = +1) WRONG RDF",
    "?",
    "?",
    "?",
    "?",
    "D17.7 (RD = +1) WRONG RDF",
    "D17.4 (RD = +1) WRONG RDF",
    "?",
    "D17.0 (RD = +1) WRONG RDF",
    "D17.2 (RD = -1)",
    "D17.6 (RD = -1)",
    "D17.7 (RD = -1)",
    "?",
    "D17.1 (RD = -1)",
    "D17.5 (RD = -1)",
    "D17.0 (RD = -1)",
    "D17.3 (RD = -1)",
    "D17.4 (RD = -1)",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "D16.2 (RD = +1) WRONG RDF",
    "D16.6 (RD = +1) WRONG RDF",
    "?",
    "?",
    "D16.1 (RD = +1) WRONG RDF",
    "D16.5 (RD = +1) WRONG RDF",
    "?",
    "D16.3 (RD = +1) WRONG RDF",
    "?",
    "?",
    "?",
    "?",
    "D09.7 (RD = +1) WRONG RDF",
    "D09.4 (RD = +1) WRONG RDF",
    "?",
    "D09.0 (RD = +1) WRONG RDF",
    "D09.2 (RD = -1)",
    "D09.6 (RD = -1)",
    "?",
    "?",
    "D09.1 (RD = -1)",
    "D09.5 (RD = -1)",
    "D09.0 (RD = -1)",
    "D09.3 (RD = -1)",
    "D09.4 (RD = -1)",
    "D09.7 (RD = -1)",
    "?",
    "?",
    "D25.7 (RD = +1) WRONG RDF",
    "D25.4 (RD = +1) WRONG RDF",
    "?",
    "D25.0 (RD = +1) WRONG RDF",
    "D25.2 (RD = -1)",
    "D25.6 (RD = -1)",
    "?",
    "?",
    "D25.1 (RD = -1)",
    "D25.5 (RD = -1)",
    "D25.0 (RD = -1)",
    "D25.3 (RD = -1)",
    "D25.4 (RD = -1)",
    "D25.7 (RD = -1)",
    "?",
    "?",
    "D00.7 (RD = -1)",
    "D00.4 (RD = -1)",
    "D00.3 (RD = -1)",
    "D00.0 (RD = -1)",
    "D00.2 (RD = -1)",
    "D00.6 (RD = -1)",
    "?",
    "?",
    "D00.1 (RD = -1)",
    "D00.5 (RD = -1)",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "D15.2 (RD = +1) WRONG RDF",
    "D15.6 (RD = +1) WRONG RDF",
    "?",
    "?",
    "D15.1 (RD = +1) WRONG RDF",
    "D15.5 (RD = +1) WRONG RDF",
    "?",
    "D15.3 (RD = +1) WRONG RDF",
    "?",
    "?",
    "?",
    "?",
    "D05.7 (RD = +1) WRONG RDF",
    "D05.4 (RD = +1) WRONG RDF",
    "?",
    "D05.0 (RD = +1) WRONG RDF",
    "D05.2 (RD = -1)",
    "D05.6 (RD = -1)",
    "?",
    "?",
    "D05.1 (RD = -1)",
    "D05.5 (RD = -1)",
    "D05.0 (RD = -1)",
    "D05.3 (RD = -1)",
    "D05.4 (RD = -1)",
    "D05.7 (RD = -1)",
    "?",
    "?",
    "D21.7 (RD = +1) WRONG RDF",
    "D21.4 (RD = +1) WRONG RDF",
    "?",
    "D21.0 (RD = +1) WRONG RDF",
    "D21.2 (RD = -1)",
    "D21.6 (RD = -1)",
    "?",
    "?",
    "D21.1 (RD = -1)",
    "D21.5 (RD = -1)",
    "D21.0 (RD = -1)",
    "D21.3 (RD = -1)",
    "D21.4 (RD = -1)",
    "D21.7 (RD = -1)",
    "?",
    "?",
    "D31.7 (RD = -1)",
    "D31.4 (RD = -1)",
    "D31.3 (RD = -1)",
    "D31.0 (RD = -1)",
    "D31.2 (RD = -1)",
    "D31.6 (RD = -1)",
    "?",
    "?",
    "D31.1 (RD = -1)",
    "D31.5 (RD = -1)",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "D13.4 (RD = +1) WRONG RDF",
    "?",
    "D13.0 (RD = +1) WRONG RDF",
    "D13.2 (RD = -1)",
    "D13.6 (RD = -1)",
    "?",
    "D13.7 (RD = +1) WRONG RDF",
    "D13.1 (RD = -1)",
    "D13.5 (RD = -1)",
    "D13.0 (RD = -1)",
    "D13.3 (RD = -1)",
    "D13.4 (RD = -1)",
    "D13.7 (RD = -1)",
    "?",
    "?",
    "D02.7 (RD = -1)",
    "D02.4 (RD = -1)",
    "D02.3 (RD = -1)",
    "D02.0 (RD = -1)",
    "D02.2 (RD = -1)",
    "D02.6 (RD = -1)",
    "?",
    "?",
    "D02.1 (RD = -1)",
    "D02.5 (RD = -1)",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "D29.7 (RD = -1)",
    "D29.4 (RD = -1)",
    "D29.3 (RD = -1)",
    "D29.0 (RD = -1)",
    "D29.2 (RD = -1)",
    "D29.6 (RD = -1)",
    "?",
    "K29.7 (RD = -1)",
    "D29.1 (RD = -1)",
    "D29.5 (RD = -1)",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "K28.5 (RD = +1) WRONG RDF",
    "K28.1 (RD = +1) WRONG RDF",
    "?",
    "?",
    "K28.6 (RD = +1) WRONG RDF",
    "K28.2 (RD = +1) WRONG RDF",
    "?",
    "K28.3 (RD = +1) WRONG RDF",
    "?",
    "?",
    "?",
    "?",
    "D03.7 (RD = +1) WRONG RDF",
    "D03.4 (RD = +1) WRONG RDF",
    "?",
    "D03.0 (RD = +1) WRONG RDF",
    "D03.2 (RD = -1)",
    "D03.6 (RD = -1)",
    "?",
    "?",
    "D03.1 (RD = -1)",
    "D03.5 (RD = -1)",
    "D03.0 (RD = -1)",
    "D03.3 (RD = -1)",
    "D03.4 (RD = -1)",
    "D03.7 (RD = -1)",
    "?",
    "?",
    "D19.7 (RD = +1) WRONG RDF",
    "D19.4 (RD = +1) WRONG RDF",
    "?",
    "D19.0 (RD = +1) WRONG RDF",
    "D19.2 (RD = -1)",
    "D19.6 (RD = -1)",
    "?",
    "?",
    "D19.1 (RD = -1)",
    "D19.5 (RD = -1)",
    "D19.0 (RD = -1)",
    "D19.3 (RD = -1)",
    "D19.4 (RD = -1)",
    "D19.7 (RD = -1)",
    "?",
    "?",
    "D24.7 (RD = -1)",
    "D24.4 (RD = -1)",
    "D24.3 (RD = -1)",
    "D24.0 (RD = -1)",
    "D24.2 (RD = -1)",
    "D24.6 (RD = -1)",
    "?",
    "?",
    "D24.1 (RD = -1)",
    "D24.5 (RD = -1)",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "D11.4 (RD = +1) WRONG RDF",
    "?",
    "D11.0 (RD = +1) WRONG RDF",
    "D11.2 (RD = -1)",
    "D11.6 (RD = -1)",
    "?",
    "D11.7 (RD = +1) WRONG RDF",
    "D11.1 (RD = -1)",
    "D11.5 (RD = -1)",
    "D11.0 (RD = -1)",
    "D11.3 (RD = -1)",
    "D11.4 (RD = -1)",
    "D11.7 (RD = -1)",
    "?",
    "?",
    "D04.7 (RD = -1)",
    "D04.4 (RD = -1)",
    "D04.3 (RD = -1)",
    "D04.0 (RD = -1)",
    "D04.2 (RD = -1)",
    "D04.6 (RD = -1)",
    "?",
    "?",
    "D04.1 (RD = -1)",
    "D04.5 (RD = -1)",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "D27.7 (RD = -1)",
    "D27.4 (RD = -1)",
    "D27.3 (RD = -1)",
    "D27.0 (RD = -1)",
    "D27.2 (RD = -1)",
    "D27.6 (RD = -1)",
    "?",
    "K27.7 (RD = -1)",
    "D27.1 (RD = -1)",
    "D27.5 (RD = -1)",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "D07.2 (RD = -1)",
    "D07.6 (RD = -1)",
    "?",
    "?",
    "D07.1 (RD = -1)",
    "D07.5 (RD = -1)",
    "D07.0 (RD = -1)",
    "D07.3 (RD = -1)",
    "D07.4 (RD = -1)",
    "D07.7 (RD = -1)",
    "?",
    "?",
    "D08.7 (RD = -1)",
    "D08.4 (RD = -1)",
    "D08.3 (RD = -1)",
    "D08.0 (RD = -1)",
    "D08.2 (RD = -1)",
    "D08.6 (RD = -1)",
    "?",
    "?",
    "D08.1 (RD = -1)",
    "D08.5 (RD = -1)",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "D23.7 (RD = -1)",
    "D23.4 (RD = -1)",
    "D23.3 (RD = -1)",
    "D23.0 (RD = -1)",
    "D23.2 (RD = -1)",
    "D23.6 (RD = -1)",
    "?",
    "K23.7 (RD = -1)",
    "D23.1 (RD = -1)",
    "D23.5 (RD = -1)",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "D23.2 (RD = +1)",
    "D23.6 (RD = +1)",
    "K23.7 (RD = +1)",
    "?",
    "D23.1 (RD = +1)",
    "D23.5 (RD = +1)",
    "D23.0 (RD = +1)",
    "D23.3 (RD = +1)",
    "D23.4 (RD = +1)",
    "D23.7 (RD = +1)",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "D08.2 (RD = +1)",
    "D08.6 (RD = +1)",
    "?",
    "?",
    "D08.1 (RD = +1)",
    "D08.5 (RD = +1)",
    "D08.0 (RD = +1)",
    "D08.3 (RD = +1)",
    "D08.4 (RD = +1)",
    "D08.7 (RD = +1)",
    "?",
    "?",
    "D07.7 (RD = +1)",
    "D07.4 (RD = +1)",
    "D07.3 (RD = +1)",
    "D07.0 (RD = +1)",
    "D07.2 (RD = +1)",
    "D07.6 (RD = +1)",
    "?",
    "?",
    "D07.1 (RD = +1)",
    "D07.5 (RD = +1)",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "D27.2 (RD = +1)",
    "D27.6 (RD = +1)",
    "K27.7 (RD = +1)",
    "?",
    "D27.1 (RD = +1)",
    "D27.5 (RD = +1)",
    "D27.0 (RD = +1)",
    "D27.3 (RD = +1)",
    "D27.4 (RD = +1)",
    "D27.7 (RD = +1)",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "D04.2 (RD = +1)",
    "D04.6 (RD = +1)",
    "?",
    "?",
    "D04.1 (RD = +1)",
    "D04.5 (RD = +1)",
    "D04.0 (RD = +1)",
    "D04.3 (RD = +1)",
    "D04.4 (RD = +1)",
    "D04.7 (RD = +1)",
    "?",
    "?",
    "D20.7 (RD = +1)",
    "D20.4 (RD = +1)",
    "D20.3 (RD = +1)",
    "D20.0 (RD = +1)",
    "D20.2 (RD = +1)",
    "D20.6 (RD = +1)",
    "D20.7 (RD = -1) WRONG RDF",
    "?",
    "D20.1 (RD = +1)",
    "D20.5 (RD = +1)",
    "D20.0 (RD = -1) WRONG RDF",
    "?",
    "D20.4 (RD = -1) WRONG RDF",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "D24.2 (RD = +1)",
    "D24.6 (RD = +1)",
    "?",
    "?",
    "D24.1 (RD = +1)",
    "D24.5 (RD = +1)",
    "D24.0 (RD = +1)",
    "D24.3 (RD = +1)",
    "D24.4 (RD = +1)",
    "D24.7 (RD = +1)",
    "?",
    "?",
    "D12.7 (RD = +1)",
    "D12.4 (RD = +1)",
    "D12.3 (RD = +1)",
    "D12.0 (RD = +1)",
    "D12.2 (RD = +1)",
    "D12.6 (RD = +1)",
    "?",
    "?",
    "D12.1 (RD = +1)",
    "D12.5 (RD = +1)",
    "D12.0 (RD = -1) WRONG RDF",
    "?",
    "D12.4 (RD = -1) WRONG RDF",
    "D12.7 (RD = -1) WRONG RDF",
    "?",
    "?",
    "D28.7 (RD = +1)",
    "D28.4 (RD = +1)",
    "D28.3 (RD = +1)",
    "D28.0 (RD = +1)",
    "D28.2 (RD = +1)",
    "D28.6 (RD = +1)",
    "?",
    "?",
    "D28.1 (RD = +1)",
    "D28.5 (RD = +1)",
    "D28.0 (RD = -1) WRONG RDF",
    "?",
    "D28.4 (RD = -1) WRONG RDF",
    "D28.7 (RD = -1) WRONG RDF",
    "?",
    "?",
    "?",
    "?",
    "K28.3 (RD = -1) WRONG RDF",
    "?",
    "K28.2 (RD = -1) WRONG RDF",
    "K28.6 (RD = -1) WRONG RDF",
    "?",
    "?",
    "K28.1 (RD = -1) WRONG RDF",
    "K28.5 (RD = -1) WRONG RDF",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "D29.2 (RD = +1)",
    "D29.6 (RD = +1)",
    "K29.7 (RD = +1)",
    "?",
    "D29.1 (RD = +1)",
    "D29.5 (RD = +1)",
    "D29.0 (RD = +1)",
    "D29.3 (RD = +1)",
    "D29.4 (RD = +1)",
    "D29.7 (RD = +1)",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "D02.2 (RD = +1)",
    "D02.6 (RD = +1)",
    "?",
    "?",
    "D02.1 (RD = +1)",
    "D02.5 (RD = +1)",
    "D02.0 (RD = +1)",
    "D02.3 (RD = +1)",
    "D02.4 (RD = +1)",
    "D02.7 (RD = +1)",
    "?",
    "?",
    "D18.7 (RD = +1)",
    "D18.4 (RD = +1)",
    "D18.3 (RD = +1)",
    "D18.0 (RD = +1)",
    "D18.2 (RD = +1)",
    "D18.6 (RD = +1)",
    "D18.7 (RD = -1) WRONG RDF",
    "?",
    "D18.1 (RD = +1)",
    "D18.5 (RD = +1)",
    "D18.0 (RD = -1) WRONG RDF",
    "?",
    "D18.4 (RD = -1) WRONG RDF",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "D31.2 (RD = +1)",
    "D31.6 (RD = +1)",
    "?",
    "?",
    "D31.1 (RD = +1)",
    "D31.5 (RD = +1)",
    "D31.0 (RD = +1)",
    "D31.3 (RD = +1)",
    "D31.4 (RD = +1)",
    "D31.7 (RD = +1)",
    "?",
    "?",
    "D10.7 (RD = +1)",
    "D10.4 (RD = +1)",
    "D10.3 (RD = +1)",
    "D10.0 (RD = +1)",
    "D10.2 (RD = +1)",
    "D10.6 (RD = +1)",
    "?",
    "?",
    "D10.1 (RD = +1)",
    "D10.5 (RD = +1)",
    "D10.0 (RD = -1) WRONG RDF",
    "?",
    "D10.4 (RD = -1) WRONG RDF",
    "D10.7 (RD = -1) WRONG RDF",
    "?",
    "?",
    "D26.7 (RD = +1)",
    "D26.4 (RD = +1)",
    "D26.3 (RD = +1)",
    "D26.0 (RD = +1)",
    "D26.2 (RD = +1)",
    "D26.6 (RD = +1)",
    "?",
    "?",
    "D26.1 (RD = +1)",
    "D26.5 (RD = +1)",
    "D26.0 (RD = -1) WRONG RDF",
    "?",
    "D26.4 (RD = -1) WRONG RDF",
    "D26.7 (RD = -1) WRONG RDF",
    "?",
    "?",
    "?",
    "?",
    "D15.3 (RD = -1) WRONG RDF",
    "?",
    "D15.2 (RD = -1) WRONG RDF",
    "D15.6 (RD = -1) WRONG RDF",
    "?",
    "?",
    "D15.1 (RD = -1) WRONG RDF",
    "D15.5 (RD = -1) WRONG RDF",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "D00.2 (RD = +1)",
    "D00.6 (RD = +1)",
    "?",
    "?",
    "D00.1 (RD = +1)",
    "D00.5 (RD = +1)",
    "D00.0 (RD = +1)",
    "D00.3 (RD = +1)",
    "D00.4 (RD = +1)",
    "D00.7 (RD = +1)",
    "?",
    "?",
    "D06.7 (RD = +1)",
    "D06.4 (RD = +1)",
    "D06.3 (RD = +1)",
    "D06.0 (RD = +1)",
    "D06.2 (RD = +1)",
    "D06.6 (RD = +1)",
    "?",
    "?",
    "D06.1 (RD = +1)",
    "D06.5 (RD = +1)",
    "D06.0 (RD = -1) WRONG RDF",
    "?",
    "D06.4 (RD = -1) WRONG RDF",
    "D06.7 (RD = -1) WRONG RDF",
    "?",
    "?",
    "D22.7 (RD = +1)",
    "D22.4 (RD = +1)",
    "D22.3 (RD = +1)",
    "D22.0 (RD = +1)",
    "D22.2 (RD = +1)",
    "D22.6 (RD = +1)",
    "?",
    "?",
    "D22.1 (RD = +1)",
    "D22.5 (RD = +1)",
    "D22.0 (RD = -1) WRONG RDF",
    "?",
    "D22.4 (RD = -1) WRONG RDF",
    "D22.7 (RD = -1) WRONG RDF",
    "?",
    "?",
    "?",
    "?",
    "D16.3 (RD = -1) WRONG RDF",
    "?",
    "D16.2 (RD = -1) WRONG RDF",
    "D16.6 (RD = -1) WRONG RDF",
    "?",
    "?",
    "D16.1 (RD = -1) WRONG RDF",
    "D16.5 (RD = -1) WRONG RDF",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "D14.4 (RD = +1)",
    "D14.3 (RD = +1)",
    "D14.0 (RD = +1)",
    "D14.2 (RD = +1)",
    "D14.6 (RD = +1)",
    "?",
    "D14.7 (RD = +1)",
    "D14.1 (RD = +1)",
    "D14.5 (RD = +1)",
    "D14.0 (RD = -1) WRONG RDF",
    "?",
    "D14.4 (RD = -1) WRONG RDF",
    "D14.7 (RD = -1) WRONG RDF",
    "?",
    "?",
    "?",
    "?",
    "D01.3 (RD = -1) WRONG RDF",
    "?",
    "D01.2 (RD = -1) WRONG RDF",
    "D01.6 (RD = -1) WRONG RDF",
    "?",
    "?",
    "D01.1 (RD = -1) WRONG RDF",
    "D01.5 (RD = -1) WRONG RDF",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "D30.3 (RD = -1) WRONG RDF",
    "?",
    "D30.2 (RD = -1) WRONG RDF",
    "D30.6 (RD = -1) WRONG RDF",
    "?",
    "?",
    "D30.1 (RD = -1) WRONG RDF",
    "D30.5 (RD = -1) WRONG RDF",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "D30.2 (RD = +1)",
    "D30.6 (RD = +1)",
    "K30.7 (RD = +1)",
    "?",
    "D30.1 (RD = +1)",
    "D30.5 (RD = +1)",
    "D30.0 (RD = +1)",
    "D30.3 (RD = +1)",
    "D30.4 (RD = +1)",
    "D30.7 (RD = +1)",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "D01.2 (RD = +1)",
    "D01.6 (RD = +1)",
    "?",
    "?",
    "D01.1 (RD = +1)",
    "D01.5 (RD = +1)",
    "D01.0 (RD = +1)",
    "D01.3 (RD = +1)",
    "D01.4 (RD = +1)",
    "D01.7 (RD = +1)",
    "?",
    "?",
    "D17.7 (RD = +1)",
    "D17.4 (RD = +1)",
    "D17.3 (RD = +1)",
    "D17.0 (RD = +1)",
    "D17.2 (RD = +1)",
    "D17.6 (RD = +1)",
    "D17.7 (RD = -1) WRONG RDF",
    "?",
    "D17.1 (RD = +1)",
    "D17.5 (RD = +1)",
    "D17.0 (RD = -1) WRONG RDF",
    "?",
    "D17.4 (RD = -1) WRONG RDF",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "D16.2 (RD = +1)",
    "D16.6 (RD = +1)",
    "?",
    "?",
    "D16.1 (RD = +1)",
    "D16.5 (RD = +1)",
    "D16.0 (RD = +1)",
    "D16.3 (RD = +1)",
    "D16.4 (RD = +1)",
    "D16.7 (RD = +1)",
    "?",
    "?",
    "D09.7 (RD = +1)",
    "D09.4 (RD = +1)",
    "D09.3 (RD = +1)",
    "D09.0 (RD = +1)",
    "D09.2 (RD = +1)",
    "D09.6 (RD = +1)",
    "?",
    "?",
    "D09.1 (RD = +1)",
    "D09.5 (RD = +1)",
    "D09.0 (RD = -1) WRONG RDF",
    "?",
    "D09.4 (RD = -1) WRONG RDF",
    "D09.7 (RD = -1) WRONG RDF",
    "?",
    "?",
    "D25.7 (RD = +1)",
    "D25.4 (RD = +1)",
    "D25.3 (RD = +1)",
    "D25.0 (RD = +1)",
    "D25.2 (RD = +1)",
    "D25.6 (RD = +1)",
    "?",
    "?",
    "D25.1 (RD = +1)",
    "D25.5 (RD = +1)",
    "D25.0 (RD = -1) WRONG RDF",
    "?",
    "D25.4 (RD = -1) WRONG RDF",
    "D25.7 (RD = -1) WRONG RDF",
    "?",
    "?",
    "?",
    "?",
    "D00.3 (RD = -1) WRONG RDF",
    "?",
    "D00.2 (RD = -1) WRONG RDF",
    "D00.6 (RD = -1) WRONG RDF",
    "?",
    "?",
    "D00.1 (RD = -1) WRONG RDF",
    "D00.5 (RD = -1) WRONG RDF",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "D15.2 (RD = +1)",
    "D15.6 (RD = +1)",
    "?",
    "?",
    "D15.1 (RD = +1)",
    "D15.5 (RD = +1)",
    "D15.0 (RD = +1)",
    "D15.3 (RD = +1)",
    "D15.4 (RD = +1)",
    "D15.7 (RD = +1)",
    "?",
    "?",
    "D05.7 (RD = +1)",
    "D05.4 (RD = +1)",
    "D05.3 (RD = +1)",
    "D05.0 (RD = +1)",
    "D05.2 (RD = +1)",
    "D05.6 (RD = +1)",
    "?",
    "?",
    "D05.1 (RD = +1)",
    "D05.5 (RD = +1)",
    "D05.0 (RD = -1) WRONG RDF",
    "?",
    "D05.4 (RD = -1) WRONG RDF",
    "D05.7 (RD = -1) WRONG RDF",
    "?",
    "?",
    "D21.7 (RD = +1)",
    "D21.4 (RD = +1)",
    "D21.3 (RD = +1)",
    "D21.0 (RD = +1)",
    "D21.2 (RD = +1)",
    "D21.6 (RD = +1)",
    "?",
    "?",
    "D21.1 (RD = +1)",
    "D21.5 (RD = +1)",
    "D21.0 (RD = -1) WRONG RDF",
    "?",
    "D21.4 (RD = -1) WRONG RDF",
    "D21.7 (RD = -1) WRONG RDF",
    "?",
    "?",
    "?",
    "?",
    "D31.3 (RD = -1) WRONG RDF",
    "?",
    "D31.2 (RD = -1) WRONG RDF",
    "D31.6 (RD = -1) WRONG RDF",
    "?",
    "?",
    "D31.1 (RD = -1) WRONG RDF",
    "D31.5 (RD = -1) WRONG RDF",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "D13.4 (RD = +1)",
    "D13.3 (RD = +1)",
    "D13.0 (RD = +1)",
    "D13.2 (RD = +1)",
    "D13.6 (RD = +1)",
    "?",
    "D13.7 (RD = +1)",
    "D13.1 (RD = +1)",
    "D13.5 (RD = +1)",
    "D13.0 (RD = -1) WRONG RDF",
    "?",
    "D13.4 (RD = -1) WRONG RDF",
    "D13.7 (RD = -1) WRONG RDF",
    "?",
    "?",
    "?",
    "?",
    "D02.3 (RD = -1) WRONG RDF",
    "?",
    "D02.2 (RD = -1) WRONG RDF",
    "D02.6 (RD = -1) WRONG RDF",
    "?",
    "?",
    "D02.1 (RD = -1) WRONG RDF",
    "D02.5 (RD = -1) WRONG RDF",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "D29.3 (RD = -1) WRONG RDF",
    "?",
    "D29.2 (RD = -1) WRONG RDF",
    "D29.6 (RD = -1) WRONG RDF",
    "?",
    "?",
    "D29.1 (RD = -1) WRONG RDF",
    "D29.5 (RD = -1) WRONG RDF",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "K28.5 (RD = +1)",
    "K28.1 (RD = +1)",
    "K28.7 (RD = +1)",
    "?",
    "K28.6 (RD = +1)",
    "K28.2 (RD = +1)",
    "K28.0 (RD = +1)",
    "K28.3 (RD = +1)",
    "K28.4 (RD = +1)",
    "?",
    "?",
    "?",
    "D03.7 (RD = +1)",
    "D03.4 (RD = +1)",
    "D03.3 (RD = +1)",
    "D03.0 (RD = +1)",
    "D03.2 (RD = +1)",
    "D03.6 (RD = +1)",
    "?",
    "?",
    "D03.1 (RD = +1)",
    "D03.5 (RD = +1)",
    "D03.0 (RD = -1) WRONG RDF",
    "?",
    "D03.4 (RD = -1) WRONG RDF",
    "D03.7 (RD = -1) WRONG RDF",
    "?",
    "?",
    "D19.7 (RD = +1)",
    "D19.4 (RD = +1)",
    "D19.3 (RD = +1)",
    "D19.0 (RD = +1)",
    "D19.2 (RD = +1)",
    "D19.6 (RD = +1)",
    "?",
    "?",
    "D19.1 (RD = +1)",
    "D19.5 (RD = +1)",
    "D19.0 (RD = -1) WRONG RDF",
    "?",
    "D19.4 (RD = -1) WRONG RDF",
    "D19.7 (RD = -1) WRONG RDF",
    "?",
    "?",
    "?",
    "?",
    "D24.3 (RD = -1) WRONG RDF",
    "?",
    "D24.2 (RD = -1) WRONG RDF",
    "D24.6 (RD = -1) WRONG RDF",
    "?",
    "?",
    "D24.1 (RD = -1) WRONG RDF",
    "D24.5 (RD = -1) WRONG RDF",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "D11.4 (RD = +1)",
    "D11.3 (RD = +1)",
    "D11.0 (RD = +1)",
    "D11.2 (RD = +1)",
    "D11.6 (RD = +1)",
    "?",
    "D11.7 (RD = +1)",
    "D11.1 (RD = +1)",
    "D11.5 (RD = +1)",
    "D11.0 (RD = -1) WRONG RDF",
    "?",
    "D11.4 (RD = -1) WRONG RDF",
    "D11.7 (RD = -1) WRONG RDF",
    "?",
    "?",
    "?",
    "?",
    "D04.3 (RD = -1) WRONG RDF",
    "?",
    "D04.2 (RD = -1) WRONG RDF",
    "D04.6 (RD = -1) WRONG RDF",
    "?",
    "?",
    "D04.1 (RD = -1) WRONG RDF",
    "D04.5 (RD = -1) WRONG RDF",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "D27.3 (RD = -1) WRONG RDF",
    "?",
    "D27.2 (RD = -1) WRONG RDF",
    "D27.6 (RD = -1) WRONG RDF",
    "?",
    "?",
    "D27.1 (RD = -1) WRONG RDF",
    "D27.5 (RD = -1) WRONG RDF",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "D07.0 (RD = -1) WRONG RDF",
    "?",
    "D07.4 (RD = -1) WRONG RDF",
    "D07.7 (RD = -1) WRONG RDF",
    "?",
    "?",
    "?",
    "?",
    "D08.3 (RD = -1) WRONG RDF",
    "?",
    "D08.2 (RD = -1) WRONG RDF",
    "D08.6 (RD = -1) WRONG RDF",
    "?",
    "?",
    "D08.1 (RD = -1) WRONG RDF",
    "D08.5 (RD = -1) WRONG RDF",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "D23.3 (RD = -1) WRONG RDF",
    "?",
    "D23.2 (RD = -1) WRONG RDF",
    "D23.6 (RD = -1) WRONG RDF",
    "?",
    "?",
    "D23.1 (RD = -1) WRONG RDF",
    "D23.5 (RD = -1) WRONG RDF",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?",
    "?"
  };

endpackage